.GLOBAL vdd! vss!


.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2

.subckt INV_X1 a zn
m_i_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
.ends INV_X1

.subckt AND2_X1 a1 a2 zn
m_i_2 net_0 a1 zn_neg vss! NMOS_VTL L=50e-9 W=210e-9
m_i_3 vss! a2 net_0 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_0 zn zn_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_5 vdd! a2 zn_neg vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_4 zn_neg a1 vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_1 zn zn_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
.ends AND2_X1

.subckt NAND2_X1 a1 a2 zn
m_i_3 zn a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_2 vdd! a1 zn vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_0 zn a1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1 net_0 a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9
.ends NAND2_X1

.subckt DEC_Read_4_13 addr[3] addr[2] addr[1] addr[0] dec_addr_bar[12] dec_addr_bar[11] dec_addr_bar[10] dec_addr_bar[9] dec_addr_bar[8] dec_addr_bar[7] dec_addr_bar[6] dec_addr_bar[5] dec_addr_bar[4] dec_addr_bar[3] dec_addr_bar[2] dec_addr_bar[1] dec_addr_bar[0]
xi3 addr[3] addr_bar[3] INV_X1
xi2 addr[2] addr_bar[2] INV_X1
xi1 addr[1] addr_bar[1] INV_X1
xi0 addr[0] addr_bar[0] INV_X1
xi11 addr[2] addr[3] net_11xx AND2_X1
xi10 addr_bar[2] addr[3] net_10xx AND2_X1
xi9 addr[2] addr_bar[3] net_01xx AND2_X1
xi8 addr_bar[2] addr_bar[3] net_00xx AND2_X1
xi7 addr[0] addr[1] net_xx11 AND2_X1
xi6 addr_bar[0] addr[1] net_xx10 AND2_X1
xi5 addr[0] addr_bar[1] net_xx01 AND2_X1
xi4 addr_bar[0] addr_bar[1] net_xx00 AND2_X1
xi24 net_xx00 net_11xx dec_addr_bar[12] NAND2_X1
xi23 net_xx11 net_10xx dec_addr_bar[11] NAND2_X1
xi22 net_xx10 net_10xx dec_addr_bar[10] NAND2_X1
xi21 net_xx01 net_10xx dec_addr_bar[9] NAND2_X1
xi20 net_xx00 net_10xx dec_addr_bar[8] NAND2_X1
xi19 net_xx11 net_01xx dec_addr_bar[7] NAND2_X1
xi18 net_xx10 net_01xx dec_addr_bar[6] NAND2_X1
xi17 net_xx01 net_01xx dec_addr_bar[5] NAND2_X1
xi16 net_xx00 net_01xx dec_addr_bar[4] NAND2_X1
xi15 net_xx11 net_00xx dec_addr_bar[3] NAND2_X1
xi14 net_xx10 net_00xx dec_addr_bar[2] NAND2_X1
xi13 net_xx01 net_00xx dec_addr_bar[1] NAND2_X1
xi12 net_xx00 net_00xx dec_addr_bar[0] NAND2_X1
.ends DEC_Read_4_13

.subckt DEC_Write_4_13 addr[3] addr[2] addr[1] addr[0] dec_addr_en[12] dec_addr_en[11] dec_addr_en[10] dec_addr_en[9] dec_addr_en[8] dec_addr_en[7] dec_addr_en[6] dec_addr_en[5] dec_addr_en[4] dec_addr_en[3] dec_addr_en[2] dec_addr_en[1] dec_addr_en[0] wr_en
xi0 addr[3] addr[2] addr[1] addr[0] dec_addr_bar[12] dec_addr_bar[11] dec_addr_bar[10] dec_addr_bar[9] dec_addr_bar[8] dec_addr_bar[7] dec_addr_bar[6] dec_addr_bar[5] dec_addr_bar[4] dec_addr_bar[3] dec_addr_bar[2] dec_addr_bar[1] dec_addr_bar[0] DEC_Read_4_13
xi1[12] dec_addr_bar[12] dec_addr[12] INV_X1
xi1[11] dec_addr_bar[11] dec_addr[11] INV_X1
xi1[10] dec_addr_bar[10] dec_addr[10] INV_X1
xi1[9] dec_addr_bar[9] dec_addr[9] INV_X1
xi1[8] dec_addr_bar[8] dec_addr[8] INV_X1
xi1[7] dec_addr_bar[7] dec_addr[7] INV_X1
xi1[6] dec_addr_bar[6] dec_addr[6] INV_X1
xi1[5] dec_addr_bar[5] dec_addr[5] INV_X1
xi1[4] dec_addr_bar[4] dec_addr[4] INV_X1
xi1[3] dec_addr_bar[3] dec_addr[3] INV_X1
xi1[2] dec_addr_bar[2] dec_addr[2] INV_X1
xi1[1] dec_addr_bar[1] dec_addr[1] INV_X1
xi1[0] dec_addr_bar[0] dec_addr[0] INV_X1
xi2[12] dec_addr[12] wr_en dec_addr_en[12] AND2_X1
xi2[11] dec_addr[11] wr_en dec_addr_en[11] AND2_X1
xi2[10] dec_addr[10] wr_en dec_addr_en[10] AND2_X1
xi2[9] dec_addr[9] wr_en dec_addr_en[9] AND2_X1
xi2[8] dec_addr[8] wr_en dec_addr_en[8] AND2_X1
xi2[7] dec_addr[7] wr_en dec_addr_en[7] AND2_X1
xi2[6] dec_addr[6] wr_en dec_addr_en[6] AND2_X1
xi2[5] dec_addr[5] wr_en dec_addr_en[5] AND2_X1
xi2[4] dec_addr[4] wr_en dec_addr_en[4] AND2_X1
xi2[3] dec_addr[3] wr_en dec_addr_en[3] AND2_X1
xi2[2] dec_addr[2] wr_en dec_addr_en[2] AND2_X1
xi2[1] dec_addr[1] wr_en dec_addr_en[1] AND2_X1
xi2[0] dec_addr[0] wr_en dec_addr_en[0] AND2_X1
.ends DEC_Write_4_13

.subckt CLKGATE_X4 ck e gck
m_i_21 vss! e net_003 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_17 net_003 net_005 net_002 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_11 net_002 net_004 net_001 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_7 net_001 net_000 vss! vss! NMOS_VTL L=50e-9 W=90e-9
m_i_45 vss! net_000 net_007b vss! NMOS_VTL L=50e-9 W=415e-9
m_i_40 net_007b ck net_006 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_40_75 net_007 ck net_006 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_45_66 vss! net_000 net_007 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_27 net_004 net_005 vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_0 vss! net_002 net_000 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_33 vss! ck net_005 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_51 gck net_006 vss! vss! NMOS_VTL L=50e-9 W=195e-9
m_i_51_7 gck net_006 vss! vss! NMOS_VTL L=50e-9 W=195e-9
m_i_51_10 gck net_006 vss! vss! NMOS_VTL L=50e-9 W=195e-9
m_i_51_7_25 gck net_006 vss! vss! NMOS_VTL L=50e-9 W=195e-9
m_i_74 net_009 net_004 net_002 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_78 vdd! e net_009 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_68 net_002 net_005 net_008 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_64 net_008 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_84 net_004 net_005 vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_57 vdd! net_002 net_000 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_90 vdd! ck net_005 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_103 vdd! net_000 net_006 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_97 net_006 ck vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_97_71 net_006 ck vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_103_74 vdd! net_000 net_006 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_109 gck net_006 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_109_4 gck net_006 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_109_24 gck net_006 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_109_4_19 gck net_006 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
.ends CLKGATE_X4

.subckt DEC_EN_4_13 ck ck_en[12] ck_en[11] ck_en[10] ck_en[9] ck_en[8] ck_en[7] ck_en[6] ck_en[5] ck_en[4] ck_en[3] ck_en[2] ck_en[1] ck_en[0] addr[3] addr[2] addr[1] addr[0] wr_en
xi0 addr[3] addr[2] addr[1] addr[0] dec_addr_en[12] dec_addr_en[11] dec_addr_en[10] dec_addr_en[9] dec_addr_en[8] dec_addr_en[7] dec_addr_en[6] dec_addr_en[5] dec_addr_en[4] dec_addr_en[3] dec_addr_en[2] dec_addr_en[1] dec_addr_en[0] wr_en DEC_Write_4_13
xi13 ck dec_addr_en[12] ck_en[12] CLKGATE_X4
xi12 ck dec_addr_en[11] ck_en[11] CLKGATE_X4
xi11 ck dec_addr_en[10] ck_en[10] CLKGATE_X4
xi10 ck dec_addr_en[9] ck_en[9] CLKGATE_X4
xi9 ck dec_addr_en[8] ck_en[8] CLKGATE_X4
xi8 ck dec_addr_en[7] ck_en[7] CLKGATE_X4
xi7 ck dec_addr_en[6] ck_en[6] CLKGATE_X4
xi6 ck dec_addr_en[5] ck_en[5] CLKGATE_X4
xi5 ck dec_addr_en[4] ck_en[4] CLKGATE_X4
xi4 ck dec_addr_en[3] ck_en[3] CLKGATE_X4
xi3 ck dec_addr_en[2] ck_en[2] CLKGATE_X4
xi2 ck dec_addr_en[1] ck_en[1] CLKGATE_X4
xi1 ck dec_addr_en[0] ck_en[0] CLKGATE_X4
.ends DEC_EN_4_13

.subckt INV_X4 a zn
m_i_0_0_x4_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_0_x4_1 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_0_x4_2 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_0_x4_3 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1_0_x4_0 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_1_0_x4_1 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_1_0_x4_2 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_1_0_x4_3 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9
.ends INV_X4

.subckt DLL_X1 d gn q
m_i_13 net_002 d vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_18 net_003 net_000 net_002 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_24 net_004 net_001 net_003 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_29 vss! net_005 net_004 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_42 q net_003 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0 net_000 gn vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_7 vss! net_000 net_001 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_35 vss! net_003 net_005 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_67 net_003 net_001 net_006 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_62 net_006 d vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_79 vdd! net_005 net_007 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_73 net_007 net_000 net_003 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_92 q net_003 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_48 net_000 gn vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_55 vdd! net_000 net_001 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_85 vdd! net_003 net_005 vdd! PMOS_VTL L=50e-9 W=90e-9
.ends DLL_X1

.subckt TBUF_X2 a en z
m_i_0_15_63 dummy1 a y vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_14_47 vss! nen dummy1 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_15 vss! a x vss! NMOS_VTL L=50e-9 W=415e-9
m_i_17 vss! en nen vss! NMOS_VTL L=50e-9 W=210e-9
m_i_0_14 vss! en x vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_6 vss! x z vss! NMOS_VTL L=50e-9 W=355e-9
m_i_0 vss! x z vss! NMOS_VTL L=50e-9 W=355e-9
m_i_24_1 dummy0 en x vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_24_0 vdd! a dummy0 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_24_0_64 vdd! a y vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_24_3 vdd! y z vdd! PMOS_VTL L=50e-9 W=540e-9
m_i_24 vdd! y z vdd! PMOS_VTL L=50e-9 W=540e-9
m_i_24_1_48 y nen vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_42 vdd! en nen vdd! PMOS_VTL L=50e-9 W=315e-9
.ends TBUF_X2

.subckt DLH_X1 d g q
m_i_13 net_002 d vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_18 net_003 net_001 net_002 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_28 vss! net_005 net_004 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_24 net_004 net_000 net_003 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_0 vss! g net_000 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_41_11 q net_003 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_7 net_001 net_000 vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_34 vss! net_003 net_005 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_66 net_003 net_000 net_006 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_61 net_006 d vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_72 net_007 net_001 net_003 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_76 vdd! net_005 net_007 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_48 vdd! g net_000 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_89_4 q net_003 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_55 net_001 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_82 vdd! net_003 net_005 vdd! PMOS_VTL L=50e-9 W=90e-9
.ends DLH_X1

.subckt cad5_13_16_REGFILE_schematic ck ck_en[12] ck_en[11] ck_en[10] ck_en[9] ck_en[8] ck_en[7] ck_en[6] ck_en[5] ck_en[4] ck_en[3] ck_en[2] ck_en[1] ck_en[0] r0_d[12] r0_d[11] r0_d[10] r0_d[9] r0_d[8] r0_d[7] r0_d[6] r0_d[5] r0_d[4] r0_d[3] r0_d[2] r0_d[1] r0_d[0] r1_d[12] r1_d[11] r1_d[10] r1_d[9] r1_d[8] r1_d[7] r1_d[6] r1_d[5] r1_d[4] r1_d[3] r1_d[2] r1_d[1] r1_d[0] rd_data_0[15] rd_data_0[14] rd_data_0[13] rd_data_0[12] rd_data_0[11] rd_data_0[10] rd_data_0[9] rd_data_0[8] rd_data_0[7] rd_data_0[6] rd_data_0[5] rd_data_0[4] rd_data_0[3] rd_data_0[2] rd_data_0[1] rd_data_0[0] rd_data_1[15] rd_data_1[14] rd_data_1[13] rd_data_1[12] rd_data_1[11] rd_data_1[10] rd_data_1[9] rd_data_1[8] rd_data_1[7] rd_data_1[6] rd_data_1[5] rd_data_1[4] rd_data_1[3] rd_data_1[2] rd_data_1[1] rd_data_1[0] wr_data[15] wr_data[14] wr_data[13] wr_data[12] wr_data[11] wr_data[10] wr_data[9] wr_data[8] wr_data[7] wr_data[6] wr_data[5] wr_data[4] wr_data[3] wr_data[2] wr_data[1] wr_data[0]
xi12[15] wr_data_preinv[15] wr_data_b[15] INV_X4
xi12[14] wr_data_preinv[14] wr_data_b[14] INV_X4
xi12[13] wr_data_preinv[13] wr_data_b[13] INV_X4
xi12[12] wr_data_preinv[12] wr_data_b[12] INV_X4
xi12[11] wr_data_preinv[11] wr_data_b[11] INV_X4
xi12[10] wr_data_preinv[10] wr_data_b[10] INV_X4
xi12[9] wr_data_preinv[9] wr_data_b[9] INV_X4
xi12[8] wr_data_preinv[8] wr_data_b[8] INV_X4
xi12[7] wr_data_preinv[7] wr_data_b[7] INV_X4
xi12[6] wr_data_preinv[6] wr_data_b[6] INV_X4
xi12[5] wr_data_preinv[5] wr_data_b[5] INV_X4
xi12[4] wr_data_preinv[4] wr_data_b[4] INV_X4
xi12[3] wr_data_preinv[3] wr_data_b[3] INV_X4
xi12[2] wr_data_preinv[2] wr_data_b[2] INV_X4
xi12[1] wr_data_preinv[1] wr_data_b[1] INV_X4
xi12[0] wr_data_preinv[0] wr_data_b[0] INV_X4
xi11[15] wr_data_prebuff[15] wr_data_preinv[15] INV_X1
xi11[14] wr_data_prebuff[14] wr_data_preinv[14] INV_X1
xi11[13] wr_data_prebuff[13] wr_data_preinv[13] INV_X1
xi11[12] wr_data_prebuff[12] wr_data_preinv[12] INV_X1
xi11[11] wr_data_prebuff[11] wr_data_preinv[11] INV_X1
xi11[10] wr_data_prebuff[10] wr_data_preinv[10] INV_X1
xi11[9] wr_data_prebuff[9] wr_data_preinv[9] INV_X1
xi11[8] wr_data_prebuff[8] wr_data_preinv[8] INV_X1
xi11[7] wr_data_prebuff[7] wr_data_preinv[7] INV_X1
xi11[6] wr_data_prebuff[6] wr_data_preinv[6] INV_X1
xi11[5] wr_data_prebuff[5] wr_data_preinv[5] INV_X1
xi11[4] wr_data_prebuff[4] wr_data_preinv[4] INV_X1
xi11[3] wr_data_prebuff[3] wr_data_preinv[3] INV_X1
xi11[2] wr_data_prebuff[2] wr_data_preinv[2] INV_X1
xi11[1] wr_data_prebuff[1] wr_data_preinv[1] INV_X1
xi11[0] wr_data_prebuff[0] wr_data_preinv[0] INV_X1
xi6[15] wr_data[15] ck wr_data_prebuff[15] DLL_X1
xi6[14] wr_data[14] ck wr_data_prebuff[14] DLL_X1
xi6[13] wr_data[13] ck wr_data_prebuff[13] DLL_X1
xi6[12] wr_data[12] ck wr_data_prebuff[12] DLL_X1
xi6[11] wr_data[11] ck wr_data_prebuff[11] DLL_X1
xi6[10] wr_data[10] ck wr_data_prebuff[10] DLL_X1
xi6[9] wr_data[9] ck wr_data_prebuff[9] DLL_X1
xi6[8] wr_data[8] ck wr_data_prebuff[8] DLL_X1
xi6[7] wr_data[7] ck wr_data_prebuff[7] DLL_X1
xi6[6] wr_data[6] ck wr_data_prebuff[6] DLL_X1
xi6[5] wr_data[5] ck wr_data_prebuff[5] DLL_X1
xi6[4] wr_data[4] ck wr_data_prebuff[4] DLL_X1
xi6[3] wr_data[3] ck wr_data_prebuff[3] DLL_X1
xi6[2] wr_data[2] ck wr_data_prebuff[2] DLL_X1
xi6[1] wr_data[1] ck wr_data_prebuff[1] DLL_X1
xi6[0] wr_data[0] ck wr_data_prebuff[0] DLL_X1
xi45[15] reg_data_10[15] r0_d[10] rd_data_0[15] TBUF_X2
xi45[14] reg_data_10[14] r0_d[10] rd_data_0[14] TBUF_X2
xi45[13] reg_data_10[13] r0_d[10] rd_data_0[13] TBUF_X2
xi45[12] reg_data_10[12] r0_d[10] rd_data_0[12] TBUF_X2
xi45[11] reg_data_10[11] r0_d[10] rd_data_0[11] TBUF_X2
xi45[10] reg_data_10[10] r0_d[10] rd_data_0[10] TBUF_X2
xi45[9] reg_data_10[9] r0_d[10] rd_data_0[9] TBUF_X2
xi45[8] reg_data_10[8] r0_d[10] rd_data_0[8] TBUF_X2
xi45[7] reg_data_10[7] r0_d[10] rd_data_0[7] TBUF_X2
xi45[6] reg_data_10[6] r0_d[10] rd_data_0[6] TBUF_X2
xi45[5] reg_data_10[5] r0_d[10] rd_data_0[5] TBUF_X2
xi45[4] reg_data_10[4] r0_d[10] rd_data_0[4] TBUF_X2
xi45[3] reg_data_10[3] r0_d[10] rd_data_0[3] TBUF_X2
xi45[2] reg_data_10[2] r0_d[10] rd_data_0[2] TBUF_X2
xi45[1] reg_data_10[1] r0_d[10] rd_data_0[1] TBUF_X2
xi45[0] reg_data_10[0] r0_d[10] rd_data_0[0] TBUF_X2
xi44[15] reg_data_10[15] r1_d[10] rd_data_1[15] TBUF_X2
xi44[14] reg_data_10[14] r1_d[10] rd_data_1[14] TBUF_X2
xi44[13] reg_data_10[13] r1_d[10] rd_data_1[13] TBUF_X2
xi44[12] reg_data_10[12] r1_d[10] rd_data_1[12] TBUF_X2
xi44[11] reg_data_10[11] r1_d[10] rd_data_1[11] TBUF_X2
xi44[10] reg_data_10[10] r1_d[10] rd_data_1[10] TBUF_X2
xi44[9] reg_data_10[9] r1_d[10] rd_data_1[9] TBUF_X2
xi44[8] reg_data_10[8] r1_d[10] rd_data_1[8] TBUF_X2
xi44[7] reg_data_10[7] r1_d[10] rd_data_1[7] TBUF_X2
xi44[6] reg_data_10[6] r1_d[10] rd_data_1[6] TBUF_X2
xi44[5] reg_data_10[5] r1_d[10] rd_data_1[5] TBUF_X2
xi44[4] reg_data_10[4] r1_d[10] rd_data_1[4] TBUF_X2
xi44[3] reg_data_10[3] r1_d[10] rd_data_1[3] TBUF_X2
xi44[2] reg_data_10[2] r1_d[10] rd_data_1[2] TBUF_X2
xi44[1] reg_data_10[1] r1_d[10] rd_data_1[1] TBUF_X2
xi44[0] reg_data_10[0] r1_d[10] rd_data_1[0] TBUF_X2
xi43[15] reg_data_11[15] r0_d[11] rd_data_0[15] TBUF_X2
xi43[14] reg_data_11[14] r0_d[11] rd_data_0[14] TBUF_X2
xi43[13] reg_data_11[13] r0_d[11] rd_data_0[13] TBUF_X2
xi43[12] reg_data_11[12] r0_d[11] rd_data_0[12] TBUF_X2
xi43[11] reg_data_11[11] r0_d[11] rd_data_0[11] TBUF_X2
xi43[10] reg_data_11[10] r0_d[11] rd_data_0[10] TBUF_X2
xi43[9] reg_data_11[9] r0_d[11] rd_data_0[9] TBUF_X2
xi43[8] reg_data_11[8] r0_d[11] rd_data_0[8] TBUF_X2
xi43[7] reg_data_11[7] r0_d[11] rd_data_0[7] TBUF_X2
xi43[6] reg_data_11[6] r0_d[11] rd_data_0[6] TBUF_X2
xi43[5] reg_data_11[5] r0_d[11] rd_data_0[5] TBUF_X2
xi43[4] reg_data_11[4] r0_d[11] rd_data_0[4] TBUF_X2
xi43[3] reg_data_11[3] r0_d[11] rd_data_0[3] TBUF_X2
xi43[2] reg_data_11[2] r0_d[11] rd_data_0[2] TBUF_X2
xi43[1] reg_data_11[1] r0_d[11] rd_data_0[1] TBUF_X2
xi43[0] reg_data_11[0] r0_d[11] rd_data_0[0] TBUF_X2
xi42[15] reg_data_11[15] r1_d[11] rd_data_1[15] TBUF_X2
xi42[14] reg_data_11[14] r1_d[11] rd_data_1[14] TBUF_X2
xi42[13] reg_data_11[13] r1_d[11] rd_data_1[13] TBUF_X2
xi42[12] reg_data_11[12] r1_d[11] rd_data_1[12] TBUF_X2
xi42[11] reg_data_11[11] r1_d[11] rd_data_1[11] TBUF_X2
xi42[10] reg_data_11[10] r1_d[11] rd_data_1[10] TBUF_X2
xi42[9] reg_data_11[9] r1_d[11] rd_data_1[9] TBUF_X2
xi42[8] reg_data_11[8] r1_d[11] rd_data_1[8] TBUF_X2
xi42[7] reg_data_11[7] r1_d[11] rd_data_1[7] TBUF_X2
xi42[6] reg_data_11[6] r1_d[11] rd_data_1[6] TBUF_X2
xi42[5] reg_data_11[5] r1_d[11] rd_data_1[5] TBUF_X2
xi42[4] reg_data_11[4] r1_d[11] rd_data_1[4] TBUF_X2
xi42[3] reg_data_11[3] r1_d[11] rd_data_1[3] TBUF_X2
xi42[2] reg_data_11[2] r1_d[11] rd_data_1[2] TBUF_X2
xi42[1] reg_data_11[1] r1_d[11] rd_data_1[1] TBUF_X2
xi42[0] reg_data_11[0] r1_d[11] rd_data_1[0] TBUF_X2
xi41[15] reg_data_12[15] r1_d[12] rd_data_1[15] TBUF_X2
xi41[14] reg_data_12[14] r1_d[12] rd_data_1[14] TBUF_X2
xi41[13] reg_data_12[13] r1_d[12] rd_data_1[13] TBUF_X2
xi41[12] reg_data_12[12] r1_d[12] rd_data_1[12] TBUF_X2
xi41[11] reg_data_12[11] r1_d[12] rd_data_1[11] TBUF_X2
xi41[10] reg_data_12[10] r1_d[12] rd_data_1[10] TBUF_X2
xi41[9] reg_data_12[9] r1_d[12] rd_data_1[9] TBUF_X2
xi41[8] reg_data_12[8] r1_d[12] rd_data_1[8] TBUF_X2
xi41[7] reg_data_12[7] r1_d[12] rd_data_1[7] TBUF_X2
xi41[6] reg_data_12[6] r1_d[12] rd_data_1[6] TBUF_X2
xi41[5] reg_data_12[5] r1_d[12] rd_data_1[5] TBUF_X2
xi41[4] reg_data_12[4] r1_d[12] rd_data_1[4] TBUF_X2
xi41[3] reg_data_12[3] r1_d[12] rd_data_1[3] TBUF_X2
xi41[2] reg_data_12[2] r1_d[12] rd_data_1[2] TBUF_X2
xi41[1] reg_data_12[1] r1_d[12] rd_data_1[1] TBUF_X2
xi41[0] reg_data_12[0] r1_d[12] rd_data_1[0] TBUF_X2
xi40[15] reg_data_12[15] r0_d[12] rd_data_0[15] TBUF_X2
xi40[14] reg_data_12[14] r0_d[12] rd_data_0[14] TBUF_X2
xi40[13] reg_data_12[13] r0_d[12] rd_data_0[13] TBUF_X2
xi40[12] reg_data_12[12] r0_d[12] rd_data_0[12] TBUF_X2
xi40[11] reg_data_12[11] r0_d[12] rd_data_0[11] TBUF_X2
xi40[10] reg_data_12[10] r0_d[12] rd_data_0[10] TBUF_X2
xi40[9] reg_data_12[9] r0_d[12] rd_data_0[9] TBUF_X2
xi40[8] reg_data_12[8] r0_d[12] rd_data_0[8] TBUF_X2
xi40[7] reg_data_12[7] r0_d[12] rd_data_0[7] TBUF_X2
xi40[6] reg_data_12[6] r0_d[12] rd_data_0[6] TBUF_X2
xi40[5] reg_data_12[5] r0_d[12] rd_data_0[5] TBUF_X2
xi40[4] reg_data_12[4] r0_d[12] rd_data_0[4] TBUF_X2
xi40[3] reg_data_12[3] r0_d[12] rd_data_0[3] TBUF_X2
xi40[2] reg_data_12[2] r0_d[12] rd_data_0[2] TBUF_X2
xi40[1] reg_data_12[1] r0_d[12] rd_data_0[1] TBUF_X2
xi40[0] reg_data_12[0] r0_d[12] rd_data_0[0] TBUF_X2
xi39[15] reg_data_9[15] r0_d[9] rd_data_0[15] TBUF_X2
xi39[14] reg_data_9[14] r0_d[9] rd_data_0[14] TBUF_X2
xi39[13] reg_data_9[13] r0_d[9] rd_data_0[13] TBUF_X2
xi39[12] reg_data_9[12] r0_d[9] rd_data_0[12] TBUF_X2
xi39[11] reg_data_9[11] r0_d[9] rd_data_0[11] TBUF_X2
xi39[10] reg_data_9[10] r0_d[9] rd_data_0[10] TBUF_X2
xi39[9] reg_data_9[9] r0_d[9] rd_data_0[9] TBUF_X2
xi39[8] reg_data_9[8] r0_d[9] rd_data_0[8] TBUF_X2
xi39[7] reg_data_9[7] r0_d[9] rd_data_0[7] TBUF_X2
xi39[6] reg_data_9[6] r0_d[9] rd_data_0[6] TBUF_X2
xi39[5] reg_data_9[5] r0_d[9] rd_data_0[5] TBUF_X2
xi39[4] reg_data_9[4] r0_d[9] rd_data_0[4] TBUF_X2
xi39[3] reg_data_9[3] r0_d[9] rd_data_0[3] TBUF_X2
xi39[2] reg_data_9[2] r0_d[9] rd_data_0[2] TBUF_X2
xi39[1] reg_data_9[1] r0_d[9] rd_data_0[1] TBUF_X2
xi39[0] reg_data_9[0] r0_d[9] rd_data_0[0] TBUF_X2
xi38[15] reg_data_9[15] r1_d[9] rd_data_1[15] TBUF_X2
xi38[14] reg_data_9[14] r1_d[9] rd_data_1[14] TBUF_X2
xi38[13] reg_data_9[13] r1_d[9] rd_data_1[13] TBUF_X2
xi38[12] reg_data_9[12] r1_d[9] rd_data_1[12] TBUF_X2
xi38[11] reg_data_9[11] r1_d[9] rd_data_1[11] TBUF_X2
xi38[10] reg_data_9[10] r1_d[9] rd_data_1[10] TBUF_X2
xi38[9] reg_data_9[9] r1_d[9] rd_data_1[9] TBUF_X2
xi38[8] reg_data_9[8] r1_d[9] rd_data_1[8] TBUF_X2
xi38[7] reg_data_9[7] r1_d[9] rd_data_1[7] TBUF_X2
xi38[6] reg_data_9[6] r1_d[9] rd_data_1[6] TBUF_X2
xi38[5] reg_data_9[5] r1_d[9] rd_data_1[5] TBUF_X2
xi38[4] reg_data_9[4] r1_d[9] rd_data_1[4] TBUF_X2
xi38[3] reg_data_9[3] r1_d[9] rd_data_1[3] TBUF_X2
xi38[2] reg_data_9[2] r1_d[9] rd_data_1[2] TBUF_X2
xi38[1] reg_data_9[1] r1_d[9] rd_data_1[1] TBUF_X2
xi38[0] reg_data_9[0] r1_d[9] rd_data_1[0] TBUF_X2
xi37[15] reg_data_8[15] r1_d[8] rd_data_1[15] TBUF_X2
xi37[14] reg_data_8[14] r1_d[8] rd_data_1[14] TBUF_X2
xi37[13] reg_data_8[13] r1_d[8] rd_data_1[13] TBUF_X2
xi37[12] reg_data_8[12] r1_d[8] rd_data_1[12] TBUF_X2
xi37[11] reg_data_8[11] r1_d[8] rd_data_1[11] TBUF_X2
xi37[10] reg_data_8[10] r1_d[8] rd_data_1[10] TBUF_X2
xi37[9] reg_data_8[9] r1_d[8] rd_data_1[9] TBUF_X2
xi37[8] reg_data_8[8] r1_d[8] rd_data_1[8] TBUF_X2
xi37[7] reg_data_8[7] r1_d[8] rd_data_1[7] TBUF_X2
xi37[6] reg_data_8[6] r1_d[8] rd_data_1[6] TBUF_X2
xi37[5] reg_data_8[5] r1_d[8] rd_data_1[5] TBUF_X2
xi37[4] reg_data_8[4] r1_d[8] rd_data_1[4] TBUF_X2
xi37[3] reg_data_8[3] r1_d[8] rd_data_1[3] TBUF_X2
xi37[2] reg_data_8[2] r1_d[8] rd_data_1[2] TBUF_X2
xi37[1] reg_data_8[1] r1_d[8] rd_data_1[1] TBUF_X2
xi37[0] reg_data_8[0] r1_d[8] rd_data_1[0] TBUF_X2
xi36[15] reg_data_8[15] r0_d[8] rd_data_0[15] TBUF_X2
xi36[14] reg_data_8[14] r0_d[8] rd_data_0[14] TBUF_X2
xi36[13] reg_data_8[13] r0_d[8] rd_data_0[13] TBUF_X2
xi36[12] reg_data_8[12] r0_d[8] rd_data_0[12] TBUF_X2
xi36[11] reg_data_8[11] r0_d[8] rd_data_0[11] TBUF_X2
xi36[10] reg_data_8[10] r0_d[8] rd_data_0[10] TBUF_X2
xi36[9] reg_data_8[9] r0_d[8] rd_data_0[9] TBUF_X2
xi36[8] reg_data_8[8] r0_d[8] rd_data_0[8] TBUF_X2
xi36[7] reg_data_8[7] r0_d[8] rd_data_0[7] TBUF_X2
xi36[6] reg_data_8[6] r0_d[8] rd_data_0[6] TBUF_X2
xi36[5] reg_data_8[5] r0_d[8] rd_data_0[5] TBUF_X2
xi36[4] reg_data_8[4] r0_d[8] rd_data_0[4] TBUF_X2
xi36[3] reg_data_8[3] r0_d[8] rd_data_0[3] TBUF_X2
xi36[2] reg_data_8[2] r0_d[8] rd_data_0[2] TBUF_X2
xi36[1] reg_data_8[1] r0_d[8] rd_data_0[1] TBUF_X2
xi36[0] reg_data_8[0] r0_d[8] rd_data_0[0] TBUF_X2
xi35[15] reg_data_7[15] r0_d[7] rd_data_0[15] TBUF_X2
xi35[14] reg_data_7[14] r0_d[7] rd_data_0[14] TBUF_X2
xi35[13] reg_data_7[13] r0_d[7] rd_data_0[13] TBUF_X2
xi35[12] reg_data_7[12] r0_d[7] rd_data_0[12] TBUF_X2
xi35[11] reg_data_7[11] r0_d[7] rd_data_0[11] TBUF_X2
xi35[10] reg_data_7[10] r0_d[7] rd_data_0[10] TBUF_X2
xi35[9] reg_data_7[9] r0_d[7] rd_data_0[9] TBUF_X2
xi35[8] reg_data_7[8] r0_d[7] rd_data_0[8] TBUF_X2
xi35[7] reg_data_7[7] r0_d[7] rd_data_0[7] TBUF_X2
xi35[6] reg_data_7[6] r0_d[7] rd_data_0[6] TBUF_X2
xi35[5] reg_data_7[5] r0_d[7] rd_data_0[5] TBUF_X2
xi35[4] reg_data_7[4] r0_d[7] rd_data_0[4] TBUF_X2
xi35[3] reg_data_7[3] r0_d[7] rd_data_0[3] TBUF_X2
xi35[2] reg_data_7[2] r0_d[7] rd_data_0[2] TBUF_X2
xi35[1] reg_data_7[1] r0_d[7] rd_data_0[1] TBUF_X2
xi35[0] reg_data_7[0] r0_d[7] rd_data_0[0] TBUF_X2
xi34[15] reg_data_7[15] r1_d[7] rd_data_1[15] TBUF_X2
xi34[14] reg_data_7[14] r1_d[7] rd_data_1[14] TBUF_X2
xi34[13] reg_data_7[13] r1_d[7] rd_data_1[13] TBUF_X2
xi34[12] reg_data_7[12] r1_d[7] rd_data_1[12] TBUF_X2
xi34[11] reg_data_7[11] r1_d[7] rd_data_1[11] TBUF_X2
xi34[10] reg_data_7[10] r1_d[7] rd_data_1[10] TBUF_X2
xi34[9] reg_data_7[9] r1_d[7] rd_data_1[9] TBUF_X2
xi34[8] reg_data_7[8] r1_d[7] rd_data_1[8] TBUF_X2
xi34[7] reg_data_7[7] r1_d[7] rd_data_1[7] TBUF_X2
xi34[6] reg_data_7[6] r1_d[7] rd_data_1[6] TBUF_X2
xi34[5] reg_data_7[5] r1_d[7] rd_data_1[5] TBUF_X2
xi34[4] reg_data_7[4] r1_d[7] rd_data_1[4] TBUF_X2
xi34[3] reg_data_7[3] r1_d[7] rd_data_1[3] TBUF_X2
xi34[2] reg_data_7[2] r1_d[7] rd_data_1[2] TBUF_X2
xi34[1] reg_data_7[1] r1_d[7] rd_data_1[1] TBUF_X2
xi34[0] reg_data_7[0] r1_d[7] rd_data_1[0] TBUF_X2
xi33[15] reg_data_6[15] r1_d[6] rd_data_1[15] TBUF_X2
xi33[14] reg_data_6[14] r1_d[6] rd_data_1[14] TBUF_X2
xi33[13] reg_data_6[13] r1_d[6] rd_data_1[13] TBUF_X2
xi33[12] reg_data_6[12] r1_d[6] rd_data_1[12] TBUF_X2
xi33[11] reg_data_6[11] r1_d[6] rd_data_1[11] TBUF_X2
xi33[10] reg_data_6[10] r1_d[6] rd_data_1[10] TBUF_X2
xi33[9] reg_data_6[9] r1_d[6] rd_data_1[9] TBUF_X2
xi33[8] reg_data_6[8] r1_d[6] rd_data_1[8] TBUF_X2
xi33[7] reg_data_6[7] r1_d[6] rd_data_1[7] TBUF_X2
xi33[6] reg_data_6[6] r1_d[6] rd_data_1[6] TBUF_X2
xi33[5] reg_data_6[5] r1_d[6] rd_data_1[5] TBUF_X2
xi33[4] reg_data_6[4] r1_d[6] rd_data_1[4] TBUF_X2
xi33[3] reg_data_6[3] r1_d[6] rd_data_1[3] TBUF_X2
xi33[2] reg_data_6[2] r1_d[6] rd_data_1[2] TBUF_X2
xi33[1] reg_data_6[1] r1_d[6] rd_data_1[1] TBUF_X2
xi33[0] reg_data_6[0] r1_d[6] rd_data_1[0] TBUF_X2
xi32[15] reg_data_6[15] r0_d[6] rd_data_0[15] TBUF_X2
xi32[14] reg_data_6[14] r0_d[6] rd_data_0[14] TBUF_X2
xi32[13] reg_data_6[13] r0_d[6] rd_data_0[13] TBUF_X2
xi32[12] reg_data_6[12] r0_d[6] rd_data_0[12] TBUF_X2
xi32[11] reg_data_6[11] r0_d[6] rd_data_0[11] TBUF_X2
xi32[10] reg_data_6[10] r0_d[6] rd_data_0[10] TBUF_X2
xi32[9] reg_data_6[9] r0_d[6] rd_data_0[9] TBUF_X2
xi32[8] reg_data_6[8] r0_d[6] rd_data_0[8] TBUF_X2
xi32[7] reg_data_6[7] r0_d[6] rd_data_0[7] TBUF_X2
xi32[6] reg_data_6[6] r0_d[6] rd_data_0[6] TBUF_X2
xi32[5] reg_data_6[5] r0_d[6] rd_data_0[5] TBUF_X2
xi32[4] reg_data_6[4] r0_d[6] rd_data_0[4] TBUF_X2
xi32[3] reg_data_6[3] r0_d[6] rd_data_0[3] TBUF_X2
xi32[2] reg_data_6[2] r0_d[6] rd_data_0[2] TBUF_X2
xi32[1] reg_data_6[1] r0_d[6] rd_data_0[1] TBUF_X2
xi32[0] reg_data_6[0] r0_d[6] rd_data_0[0] TBUF_X2
xi31[15] reg_data_5[15] r1_d[5] rd_data_1[15] TBUF_X2
xi31[14] reg_data_5[14] r1_d[5] rd_data_1[14] TBUF_X2
xi31[13] reg_data_5[13] r1_d[5] rd_data_1[13] TBUF_X2
xi31[12] reg_data_5[12] r1_d[5] rd_data_1[12] TBUF_X2
xi31[11] reg_data_5[11] r1_d[5] rd_data_1[11] TBUF_X2
xi31[10] reg_data_5[10] r1_d[5] rd_data_1[10] TBUF_X2
xi31[9] reg_data_5[9] r1_d[5] rd_data_1[9] TBUF_X2
xi31[8] reg_data_5[8] r1_d[5] rd_data_1[8] TBUF_X2
xi31[7] reg_data_5[7] r1_d[5] rd_data_1[7] TBUF_X2
xi31[6] reg_data_5[6] r1_d[5] rd_data_1[6] TBUF_X2
xi31[5] reg_data_5[5] r1_d[5] rd_data_1[5] TBUF_X2
xi31[4] reg_data_5[4] r1_d[5] rd_data_1[4] TBUF_X2
xi31[3] reg_data_5[3] r1_d[5] rd_data_1[3] TBUF_X2
xi31[2] reg_data_5[2] r1_d[5] rd_data_1[2] TBUF_X2
xi31[1] reg_data_5[1] r1_d[5] rd_data_1[1] TBUF_X2
xi31[0] reg_data_5[0] r1_d[5] rd_data_1[0] TBUF_X2
xi30[15] reg_data_5[15] r0_d[5] rd_data_0[15] TBUF_X2
xi30[14] reg_data_5[14] r0_d[5] rd_data_0[14] TBUF_X2
xi30[13] reg_data_5[13] r0_d[5] rd_data_0[13] TBUF_X2
xi30[12] reg_data_5[12] r0_d[5] rd_data_0[12] TBUF_X2
xi30[11] reg_data_5[11] r0_d[5] rd_data_0[11] TBUF_X2
xi30[10] reg_data_5[10] r0_d[5] rd_data_0[10] TBUF_X2
xi30[9] reg_data_5[9] r0_d[5] rd_data_0[9] TBUF_X2
xi30[8] reg_data_5[8] r0_d[5] rd_data_0[8] TBUF_X2
xi30[7] reg_data_5[7] r0_d[5] rd_data_0[7] TBUF_X2
xi30[6] reg_data_5[6] r0_d[5] rd_data_0[6] TBUF_X2
xi30[5] reg_data_5[5] r0_d[5] rd_data_0[5] TBUF_X2
xi30[4] reg_data_5[4] r0_d[5] rd_data_0[4] TBUF_X2
xi30[3] reg_data_5[3] r0_d[5] rd_data_0[3] TBUF_X2
xi30[2] reg_data_5[2] r0_d[5] rd_data_0[2] TBUF_X2
xi30[1] reg_data_5[1] r0_d[5] rd_data_0[1] TBUF_X2
xi30[0] reg_data_5[0] r0_d[5] rd_data_0[0] TBUF_X2
xi29[15] reg_data_4[15] r1_d[4] rd_data_1[15] TBUF_X2
xi29[14] reg_data_4[14] r1_d[4] rd_data_1[14] TBUF_X2
xi29[13] reg_data_4[13] r1_d[4] rd_data_1[13] TBUF_X2
xi29[12] reg_data_4[12] r1_d[4] rd_data_1[12] TBUF_X2
xi29[11] reg_data_4[11] r1_d[4] rd_data_1[11] TBUF_X2
xi29[10] reg_data_4[10] r1_d[4] rd_data_1[10] TBUF_X2
xi29[9] reg_data_4[9] r1_d[4] rd_data_1[9] TBUF_X2
xi29[8] reg_data_4[8] r1_d[4] rd_data_1[8] TBUF_X2
xi29[7] reg_data_4[7] r1_d[4] rd_data_1[7] TBUF_X2
xi29[6] reg_data_4[6] r1_d[4] rd_data_1[6] TBUF_X2
xi29[5] reg_data_4[5] r1_d[4] rd_data_1[5] TBUF_X2
xi29[4] reg_data_4[4] r1_d[4] rd_data_1[4] TBUF_X2
xi29[3] reg_data_4[3] r1_d[4] rd_data_1[3] TBUF_X2
xi29[2] reg_data_4[2] r1_d[4] rd_data_1[2] TBUF_X2
xi29[1] reg_data_4[1] r1_d[4] rd_data_1[1] TBUF_X2
xi29[0] reg_data_4[0] r1_d[4] rd_data_1[0] TBUF_X2
xi28[15] reg_data_4[15] r0_d[4] rd_data_0[15] TBUF_X2
xi28[14] reg_data_4[14] r0_d[4] rd_data_0[14] TBUF_X2
xi28[13] reg_data_4[13] r0_d[4] rd_data_0[13] TBUF_X2
xi28[12] reg_data_4[12] r0_d[4] rd_data_0[12] TBUF_X2
xi28[11] reg_data_4[11] r0_d[4] rd_data_0[11] TBUF_X2
xi28[10] reg_data_4[10] r0_d[4] rd_data_0[10] TBUF_X2
xi28[9] reg_data_4[9] r0_d[4] rd_data_0[9] TBUF_X2
xi28[8] reg_data_4[8] r0_d[4] rd_data_0[8] TBUF_X2
xi28[7] reg_data_4[7] r0_d[4] rd_data_0[7] TBUF_X2
xi28[6] reg_data_4[6] r0_d[4] rd_data_0[6] TBUF_X2
xi28[5] reg_data_4[5] r0_d[4] rd_data_0[5] TBUF_X2
xi28[4] reg_data_4[4] r0_d[4] rd_data_0[4] TBUF_X2
xi28[3] reg_data_4[3] r0_d[4] rd_data_0[3] TBUF_X2
xi28[2] reg_data_4[2] r0_d[4] rd_data_0[2] TBUF_X2
xi28[1] reg_data_4[1] r0_d[4] rd_data_0[1] TBUF_X2
xi28[0] reg_data_4[0] r0_d[4] rd_data_0[0] TBUF_X2
xi27[15] reg_data_3[15] r0_d[3] rd_data_0[15] TBUF_X2
xi27[14] reg_data_3[14] r0_d[3] rd_data_0[14] TBUF_X2
xi27[13] reg_data_3[13] r0_d[3] rd_data_0[13] TBUF_X2
xi27[12] reg_data_3[12] r0_d[3] rd_data_0[12] TBUF_X2
xi27[11] reg_data_3[11] r0_d[3] rd_data_0[11] TBUF_X2
xi27[10] reg_data_3[10] r0_d[3] rd_data_0[10] TBUF_X2
xi27[9] reg_data_3[9] r0_d[3] rd_data_0[9] TBUF_X2
xi27[8] reg_data_3[8] r0_d[3] rd_data_0[8] TBUF_X2
xi27[7] reg_data_3[7] r0_d[3] rd_data_0[7] TBUF_X2
xi27[6] reg_data_3[6] r0_d[3] rd_data_0[6] TBUF_X2
xi27[5] reg_data_3[5] r0_d[3] rd_data_0[5] TBUF_X2
xi27[4] reg_data_3[4] r0_d[3] rd_data_0[4] TBUF_X2
xi27[3] reg_data_3[3] r0_d[3] rd_data_0[3] TBUF_X2
xi27[2] reg_data_3[2] r0_d[3] rd_data_0[2] TBUF_X2
xi27[1] reg_data_3[1] r0_d[3] rd_data_0[1] TBUF_X2
xi27[0] reg_data_3[0] r0_d[3] rd_data_0[0] TBUF_X2
xi26[15] reg_data_3[15] r1_d[3] rd_data_1[15] TBUF_X2
xi26[14] reg_data_3[14] r1_d[3] rd_data_1[14] TBUF_X2
xi26[13] reg_data_3[13] r1_d[3] rd_data_1[13] TBUF_X2
xi26[12] reg_data_3[12] r1_d[3] rd_data_1[12] TBUF_X2
xi26[11] reg_data_3[11] r1_d[3] rd_data_1[11] TBUF_X2
xi26[10] reg_data_3[10] r1_d[3] rd_data_1[10] TBUF_X2
xi26[9] reg_data_3[9] r1_d[3] rd_data_1[9] TBUF_X2
xi26[8] reg_data_3[8] r1_d[3] rd_data_1[8] TBUF_X2
xi26[7] reg_data_3[7] r1_d[3] rd_data_1[7] TBUF_X2
xi26[6] reg_data_3[6] r1_d[3] rd_data_1[6] TBUF_X2
xi26[5] reg_data_3[5] r1_d[3] rd_data_1[5] TBUF_X2
xi26[4] reg_data_3[4] r1_d[3] rd_data_1[4] TBUF_X2
xi26[3] reg_data_3[3] r1_d[3] rd_data_1[3] TBUF_X2
xi26[2] reg_data_3[2] r1_d[3] rd_data_1[2] TBUF_X2
xi26[1] reg_data_3[1] r1_d[3] rd_data_1[1] TBUF_X2
xi26[0] reg_data_3[0] r1_d[3] rd_data_1[0] TBUF_X2
xi25[15] reg_data_2[15] r1_d[2] rd_data_1[15] TBUF_X2
xi25[14] reg_data_2[14] r1_d[2] rd_data_1[14] TBUF_X2
xi25[13] reg_data_2[13] r1_d[2] rd_data_1[13] TBUF_X2
xi25[12] reg_data_2[12] r1_d[2] rd_data_1[12] TBUF_X2
xi25[11] reg_data_2[11] r1_d[2] rd_data_1[11] TBUF_X2
xi25[10] reg_data_2[10] r1_d[2] rd_data_1[10] TBUF_X2
xi25[9] reg_data_2[9] r1_d[2] rd_data_1[9] TBUF_X2
xi25[8] reg_data_2[8] r1_d[2] rd_data_1[8] TBUF_X2
xi25[7] reg_data_2[7] r1_d[2] rd_data_1[7] TBUF_X2
xi25[6] reg_data_2[6] r1_d[2] rd_data_1[6] TBUF_X2
xi25[5] reg_data_2[5] r1_d[2] rd_data_1[5] TBUF_X2
xi25[4] reg_data_2[4] r1_d[2] rd_data_1[4] TBUF_X2
xi25[3] reg_data_2[3] r1_d[2] rd_data_1[3] TBUF_X2
xi25[2] reg_data_2[2] r1_d[2] rd_data_1[2] TBUF_X2
xi25[1] reg_data_2[1] r1_d[2] rd_data_1[1] TBUF_X2
xi25[0] reg_data_2[0] r1_d[2] rd_data_1[0] TBUF_X2
xi3[15] reg_data_0[15] r1_d[0] rd_data_1[15] TBUF_X2
xi3[14] reg_data_0[14] r1_d[0] rd_data_1[14] TBUF_X2
xi3[13] reg_data_0[13] r1_d[0] rd_data_1[13] TBUF_X2
xi3[12] reg_data_0[12] r1_d[0] rd_data_1[12] TBUF_X2
xi3[11] reg_data_0[11] r1_d[0] rd_data_1[11] TBUF_X2
xi3[10] reg_data_0[10] r1_d[0] rd_data_1[10] TBUF_X2
xi3[9] reg_data_0[9] r1_d[0] rd_data_1[9] TBUF_X2
xi3[8] reg_data_0[8] r1_d[0] rd_data_1[8] TBUF_X2
xi3[7] reg_data_0[7] r1_d[0] rd_data_1[7] TBUF_X2
xi3[6] reg_data_0[6] r1_d[0] rd_data_1[6] TBUF_X2
xi3[5] reg_data_0[5] r1_d[0] rd_data_1[5] TBUF_X2
xi3[4] reg_data_0[4] r1_d[0] rd_data_1[4] TBUF_X2
xi3[3] reg_data_0[3] r1_d[0] rd_data_1[3] TBUF_X2
xi3[2] reg_data_0[2] r1_d[0] rd_data_1[2] TBUF_X2
xi3[1] reg_data_0[1] r1_d[0] rd_data_1[1] TBUF_X2
xi3[0] reg_data_0[0] r1_d[0] rd_data_1[0] TBUF_X2
xi24[15] reg_data_2[15] r0_d[2] rd_data_0[15] TBUF_X2
xi24[14] reg_data_2[14] r0_d[2] rd_data_0[14] TBUF_X2
xi24[13] reg_data_2[13] r0_d[2] rd_data_0[13] TBUF_X2
xi24[12] reg_data_2[12] r0_d[2] rd_data_0[12] TBUF_X2
xi24[11] reg_data_2[11] r0_d[2] rd_data_0[11] TBUF_X2
xi24[10] reg_data_2[10] r0_d[2] rd_data_0[10] TBUF_X2
xi24[9] reg_data_2[9] r0_d[2] rd_data_0[9] TBUF_X2
xi24[8] reg_data_2[8] r0_d[2] rd_data_0[8] TBUF_X2
xi24[7] reg_data_2[7] r0_d[2] rd_data_0[7] TBUF_X2
xi24[6] reg_data_2[6] r0_d[2] rd_data_0[6] TBUF_X2
xi24[5] reg_data_2[5] r0_d[2] rd_data_0[5] TBUF_X2
xi24[4] reg_data_2[4] r0_d[2] rd_data_0[4] TBUF_X2
xi24[3] reg_data_2[3] r0_d[2] rd_data_0[3] TBUF_X2
xi24[2] reg_data_2[2] r0_d[2] rd_data_0[2] TBUF_X2
xi24[1] reg_data_2[1] r0_d[2] rd_data_0[1] TBUF_X2
xi24[0] reg_data_2[0] r0_d[2] rd_data_0[0] TBUF_X2
xi4[15] reg_data_0[15] r0_d[0] rd_data_0[15] TBUF_X2
xi4[14] reg_data_0[14] r0_d[0] rd_data_0[14] TBUF_X2
xi4[13] reg_data_0[13] r0_d[0] rd_data_0[13] TBUF_X2
xi4[12] reg_data_0[12] r0_d[0] rd_data_0[12] TBUF_X2
xi4[11] reg_data_0[11] r0_d[0] rd_data_0[11] TBUF_X2
xi4[10] reg_data_0[10] r0_d[0] rd_data_0[10] TBUF_X2
xi4[9] reg_data_0[9] r0_d[0] rd_data_0[9] TBUF_X2
xi4[8] reg_data_0[8] r0_d[0] rd_data_0[8] TBUF_X2
xi4[7] reg_data_0[7] r0_d[0] rd_data_0[7] TBUF_X2
xi4[6] reg_data_0[6] r0_d[0] rd_data_0[6] TBUF_X2
xi4[5] reg_data_0[5] r0_d[0] rd_data_0[5] TBUF_X2
xi4[4] reg_data_0[4] r0_d[0] rd_data_0[4] TBUF_X2
xi4[3] reg_data_0[3] r0_d[0] rd_data_0[3] TBUF_X2
xi4[2] reg_data_0[2] r0_d[0] rd_data_0[2] TBUF_X2
xi4[1] reg_data_0[1] r0_d[0] rd_data_0[1] TBUF_X2
xi4[0] reg_data_0[0] r0_d[0] rd_data_0[0] TBUF_X2
xi10[15] reg_data_1[15] r1_d[1] rd_data_1[15] TBUF_X2
xi10[14] reg_data_1[14] r1_d[1] rd_data_1[14] TBUF_X2
xi10[13] reg_data_1[13] r1_d[1] rd_data_1[13] TBUF_X2
xi10[12] reg_data_1[12] r1_d[1] rd_data_1[12] TBUF_X2
xi10[11] reg_data_1[11] r1_d[1] rd_data_1[11] TBUF_X2
xi10[10] reg_data_1[10] r1_d[1] rd_data_1[10] TBUF_X2
xi10[9] reg_data_1[9] r1_d[1] rd_data_1[9] TBUF_X2
xi10[8] reg_data_1[8] r1_d[1] rd_data_1[8] TBUF_X2
xi10[7] reg_data_1[7] r1_d[1] rd_data_1[7] TBUF_X2
xi10[6] reg_data_1[6] r1_d[1] rd_data_1[6] TBUF_X2
xi10[5] reg_data_1[5] r1_d[1] rd_data_1[5] TBUF_X2
xi10[4] reg_data_1[4] r1_d[1] rd_data_1[4] TBUF_X2
xi10[3] reg_data_1[3] r1_d[1] rd_data_1[3] TBUF_X2
xi10[2] reg_data_1[2] r1_d[1] rd_data_1[2] TBUF_X2
xi10[1] reg_data_1[1] r1_d[1] rd_data_1[1] TBUF_X2
xi10[0] reg_data_1[0] r1_d[1] rd_data_1[0] TBUF_X2
xi9[15] reg_data_1[15] r0_d[1] rd_data_0[15] TBUF_X2
xi9[14] reg_data_1[14] r0_d[1] rd_data_0[14] TBUF_X2
xi9[13] reg_data_1[13] r0_d[1] rd_data_0[13] TBUF_X2
xi9[12] reg_data_1[12] r0_d[1] rd_data_0[12] TBUF_X2
xi9[11] reg_data_1[11] r0_d[1] rd_data_0[11] TBUF_X2
xi9[10] reg_data_1[10] r0_d[1] rd_data_0[10] TBUF_X2
xi9[9] reg_data_1[9] r0_d[1] rd_data_0[9] TBUF_X2
xi9[8] reg_data_1[8] r0_d[1] rd_data_0[8] TBUF_X2
xi9[7] reg_data_1[7] r0_d[1] rd_data_0[7] TBUF_X2
xi9[6] reg_data_1[6] r0_d[1] rd_data_0[6] TBUF_X2
xi9[5] reg_data_1[5] r0_d[1] rd_data_0[5] TBUF_X2
xi9[4] reg_data_1[4] r0_d[1] rd_data_0[4] TBUF_X2
xi9[3] reg_data_1[3] r0_d[1] rd_data_0[3] TBUF_X2
xi9[2] reg_data_1[2] r0_d[1] rd_data_0[2] TBUF_X2
xi9[1] reg_data_1[1] r0_d[1] rd_data_0[1] TBUF_X2
xi9[0] reg_data_1[0] r0_d[1] rd_data_0[0] TBUF_X2
xi23[15] wr_data_b[15] ck_en[12] reg_data_12[15] DLH_X1
xi23[14] wr_data_b[14] ck_en[12] reg_data_12[14] DLH_X1
xi23[13] wr_data_b[13] ck_en[12] reg_data_12[13] DLH_X1
xi23[12] wr_data_b[12] ck_en[12] reg_data_12[12] DLH_X1
xi23[11] wr_data_b[11] ck_en[12] reg_data_12[11] DLH_X1
xi23[10] wr_data_b[10] ck_en[12] reg_data_12[10] DLH_X1
xi23[9] wr_data_b[9] ck_en[12] reg_data_12[9] DLH_X1
xi23[8] wr_data_b[8] ck_en[12] reg_data_12[8] DLH_X1
xi23[7] wr_data_b[7] ck_en[12] reg_data_12[7] DLH_X1
xi23[6] wr_data_b[6] ck_en[12] reg_data_12[6] DLH_X1
xi23[5] wr_data_b[5] ck_en[12] reg_data_12[5] DLH_X1
xi23[4] wr_data_b[4] ck_en[12] reg_data_12[4] DLH_X1
xi23[3] wr_data_b[3] ck_en[12] reg_data_12[3] DLH_X1
xi23[2] wr_data_b[2] ck_en[12] reg_data_12[2] DLH_X1
xi23[1] wr_data_b[1] ck_en[12] reg_data_12[1] DLH_X1
xi23[0] wr_data_b[0] ck_en[12] reg_data_12[0] DLH_X1
xi22[15] wr_data_b[15] ck_en[7] reg_data_7[15] DLH_X1
xi22[14] wr_data_b[14] ck_en[7] reg_data_7[14] DLH_X1
xi22[13] wr_data_b[13] ck_en[7] reg_data_7[13] DLH_X1
xi22[12] wr_data_b[12] ck_en[7] reg_data_7[12] DLH_X1
xi22[11] wr_data_b[11] ck_en[7] reg_data_7[11] DLH_X1
xi22[10] wr_data_b[10] ck_en[7] reg_data_7[10] DLH_X1
xi22[9] wr_data_b[9] ck_en[7] reg_data_7[9] DLH_X1
xi22[8] wr_data_b[8] ck_en[7] reg_data_7[8] DLH_X1
xi22[7] wr_data_b[7] ck_en[7] reg_data_7[7] DLH_X1
xi22[6] wr_data_b[6] ck_en[7] reg_data_7[6] DLH_X1
xi22[5] wr_data_b[5] ck_en[7] reg_data_7[5] DLH_X1
xi22[4] wr_data_b[4] ck_en[7] reg_data_7[4] DLH_X1
xi22[3] wr_data_b[3] ck_en[7] reg_data_7[3] DLH_X1
xi22[2] wr_data_b[2] ck_en[7] reg_data_7[2] DLH_X1
xi22[1] wr_data_b[1] ck_en[7] reg_data_7[1] DLH_X1
xi22[0] wr_data_b[0] ck_en[7] reg_data_7[0] DLH_X1
xi21[15] wr_data_b[15] ck_en[8] reg_data_8[15] DLH_X1
xi21[14] wr_data_b[14] ck_en[8] reg_data_8[14] DLH_X1
xi21[13] wr_data_b[13] ck_en[8] reg_data_8[13] DLH_X1
xi21[12] wr_data_b[12] ck_en[8] reg_data_8[12] DLH_X1
xi21[11] wr_data_b[11] ck_en[8] reg_data_8[11] DLH_X1
xi21[10] wr_data_b[10] ck_en[8] reg_data_8[10] DLH_X1
xi21[9] wr_data_b[9] ck_en[8] reg_data_8[9] DLH_X1
xi21[8] wr_data_b[8] ck_en[8] reg_data_8[8] DLH_X1
xi21[7] wr_data_b[7] ck_en[8] reg_data_8[7] DLH_X1
xi21[6] wr_data_b[6] ck_en[8] reg_data_8[6] DLH_X1
xi21[5] wr_data_b[5] ck_en[8] reg_data_8[5] DLH_X1
xi21[4] wr_data_b[4] ck_en[8] reg_data_8[4] DLH_X1
xi21[3] wr_data_b[3] ck_en[8] reg_data_8[3] DLH_X1
xi21[2] wr_data_b[2] ck_en[8] reg_data_8[2] DLH_X1
xi21[1] wr_data_b[1] ck_en[8] reg_data_8[1] DLH_X1
xi21[0] wr_data_b[0] ck_en[8] reg_data_8[0] DLH_X1
xi20[15] wr_data_b[15] ck_en[9] reg_data_9[15] DLH_X1
xi20[14] wr_data_b[14] ck_en[9] reg_data_9[14] DLH_X1
xi20[13] wr_data_b[13] ck_en[9] reg_data_9[13] DLH_X1
xi20[12] wr_data_b[12] ck_en[9] reg_data_9[12] DLH_X1
xi20[11] wr_data_b[11] ck_en[9] reg_data_9[11] DLH_X1
xi20[10] wr_data_b[10] ck_en[9] reg_data_9[10] DLH_X1
xi20[9] wr_data_b[9] ck_en[9] reg_data_9[9] DLH_X1
xi20[8] wr_data_b[8] ck_en[9] reg_data_9[8] DLH_X1
xi20[7] wr_data_b[7] ck_en[9] reg_data_9[7] DLH_X1
xi20[6] wr_data_b[6] ck_en[9] reg_data_9[6] DLH_X1
xi20[5] wr_data_b[5] ck_en[9] reg_data_9[5] DLH_X1
xi20[4] wr_data_b[4] ck_en[9] reg_data_9[4] DLH_X1
xi20[3] wr_data_b[3] ck_en[9] reg_data_9[3] DLH_X1
xi20[2] wr_data_b[2] ck_en[9] reg_data_9[2] DLH_X1
xi20[1] wr_data_b[1] ck_en[9] reg_data_9[1] DLH_X1
xi20[0] wr_data_b[0] ck_en[9] reg_data_9[0] DLH_X1
xi19[15] wr_data_b[15] ck_en[11] reg_data_11[15] DLH_X1
xi19[14] wr_data_b[14] ck_en[11] reg_data_11[14] DLH_X1
xi19[13] wr_data_b[13] ck_en[11] reg_data_11[13] DLH_X1
xi19[12] wr_data_b[12] ck_en[11] reg_data_11[12] DLH_X1
xi19[11] wr_data_b[11] ck_en[11] reg_data_11[11] DLH_X1
xi19[10] wr_data_b[10] ck_en[11] reg_data_11[10] DLH_X1
xi19[9] wr_data_b[9] ck_en[11] reg_data_11[9] DLH_X1
xi19[8] wr_data_b[8] ck_en[11] reg_data_11[8] DLH_X1
xi19[7] wr_data_b[7] ck_en[11] reg_data_11[7] DLH_X1
xi19[6] wr_data_b[6] ck_en[11] reg_data_11[6] DLH_X1
xi19[5] wr_data_b[5] ck_en[11] reg_data_11[5] DLH_X1
xi19[4] wr_data_b[4] ck_en[11] reg_data_11[4] DLH_X1
xi19[3] wr_data_b[3] ck_en[11] reg_data_11[3] DLH_X1
xi19[2] wr_data_b[2] ck_en[11] reg_data_11[2] DLH_X1
xi19[1] wr_data_b[1] ck_en[11] reg_data_11[1] DLH_X1
xi19[0] wr_data_b[0] ck_en[11] reg_data_11[0] DLH_X1
xi18[15] wr_data_b[15] ck_en[10] reg_data_10[15] DLH_X1
xi18[14] wr_data_b[14] ck_en[10] reg_data_10[14] DLH_X1
xi18[13] wr_data_b[13] ck_en[10] reg_data_10[13] DLH_X1
xi18[12] wr_data_b[12] ck_en[10] reg_data_10[12] DLH_X1
xi18[11] wr_data_b[11] ck_en[10] reg_data_10[11] DLH_X1
xi18[10] wr_data_b[10] ck_en[10] reg_data_10[10] DLH_X1
xi18[9] wr_data_b[9] ck_en[10] reg_data_10[9] DLH_X1
xi18[8] wr_data_b[8] ck_en[10] reg_data_10[8] DLH_X1
xi18[7] wr_data_b[7] ck_en[10] reg_data_10[7] DLH_X1
xi18[6] wr_data_b[6] ck_en[10] reg_data_10[6] DLH_X1
xi18[5] wr_data_b[5] ck_en[10] reg_data_10[5] DLH_X1
xi18[4] wr_data_b[4] ck_en[10] reg_data_10[4] DLH_X1
xi18[3] wr_data_b[3] ck_en[10] reg_data_10[3] DLH_X1
xi18[2] wr_data_b[2] ck_en[10] reg_data_10[2] DLH_X1
xi18[1] wr_data_b[1] ck_en[10] reg_data_10[1] DLH_X1
xi18[0] wr_data_b[0] ck_en[10] reg_data_10[0] DLH_X1
xi17[15] wr_data_b[15] ck_en[6] reg_data_6[15] DLH_X1
xi17[14] wr_data_b[14] ck_en[6] reg_data_6[14] DLH_X1
xi17[13] wr_data_b[13] ck_en[6] reg_data_6[13] DLH_X1
xi17[12] wr_data_b[12] ck_en[6] reg_data_6[12] DLH_X1
xi17[11] wr_data_b[11] ck_en[6] reg_data_6[11] DLH_X1
xi17[10] wr_data_b[10] ck_en[6] reg_data_6[10] DLH_X1
xi17[9] wr_data_b[9] ck_en[6] reg_data_6[9] DLH_X1
xi17[8] wr_data_b[8] ck_en[6] reg_data_6[8] DLH_X1
xi17[7] wr_data_b[7] ck_en[6] reg_data_6[7] DLH_X1
xi17[6] wr_data_b[6] ck_en[6] reg_data_6[6] DLH_X1
xi17[5] wr_data_b[5] ck_en[6] reg_data_6[5] DLH_X1
xi17[4] wr_data_b[4] ck_en[6] reg_data_6[4] DLH_X1
xi17[3] wr_data_b[3] ck_en[6] reg_data_6[3] DLH_X1
xi17[2] wr_data_b[2] ck_en[6] reg_data_6[2] DLH_X1
xi17[1] wr_data_b[1] ck_en[6] reg_data_6[1] DLH_X1
xi17[0] wr_data_b[0] ck_en[6] reg_data_6[0] DLH_X1
xi16[15] wr_data_b[15] ck_en[5] reg_data_5[15] DLH_X1
xi16[14] wr_data_b[14] ck_en[5] reg_data_5[14] DLH_X1
xi16[13] wr_data_b[13] ck_en[5] reg_data_5[13] DLH_X1
xi16[12] wr_data_b[12] ck_en[5] reg_data_5[12] DLH_X1
xi16[11] wr_data_b[11] ck_en[5] reg_data_5[11] DLH_X1
xi16[10] wr_data_b[10] ck_en[5] reg_data_5[10] DLH_X1
xi16[9] wr_data_b[9] ck_en[5] reg_data_5[9] DLH_X1
xi16[8] wr_data_b[8] ck_en[5] reg_data_5[8] DLH_X1
xi16[7] wr_data_b[7] ck_en[5] reg_data_5[7] DLH_X1
xi16[6] wr_data_b[6] ck_en[5] reg_data_5[6] DLH_X1
xi16[5] wr_data_b[5] ck_en[5] reg_data_5[5] DLH_X1
xi16[4] wr_data_b[4] ck_en[5] reg_data_5[4] DLH_X1
xi16[3] wr_data_b[3] ck_en[5] reg_data_5[3] DLH_X1
xi16[2] wr_data_b[2] ck_en[5] reg_data_5[2] DLH_X1
xi16[1] wr_data_b[1] ck_en[5] reg_data_5[1] DLH_X1
xi16[0] wr_data_b[0] ck_en[5] reg_data_5[0] DLH_X1
xi15[15] wr_data_b[15] ck_en[4] reg_data_4[15] DLH_X1
xi15[14] wr_data_b[14] ck_en[4] reg_data_4[14] DLH_X1
xi15[13] wr_data_b[13] ck_en[4] reg_data_4[13] DLH_X1
xi15[12] wr_data_b[12] ck_en[4] reg_data_4[12] DLH_X1
xi15[11] wr_data_b[11] ck_en[4] reg_data_4[11] DLH_X1
xi15[10] wr_data_b[10] ck_en[4] reg_data_4[10] DLH_X1
xi15[9] wr_data_b[9] ck_en[4] reg_data_4[9] DLH_X1
xi15[8] wr_data_b[8] ck_en[4] reg_data_4[8] DLH_X1
xi15[7] wr_data_b[7] ck_en[4] reg_data_4[7] DLH_X1
xi15[6] wr_data_b[6] ck_en[4] reg_data_4[6] DLH_X1
xi15[5] wr_data_b[5] ck_en[4] reg_data_4[5] DLH_X1
xi15[4] wr_data_b[4] ck_en[4] reg_data_4[4] DLH_X1
xi15[3] wr_data_b[3] ck_en[4] reg_data_4[3] DLH_X1
xi15[2] wr_data_b[2] ck_en[4] reg_data_4[2] DLH_X1
xi15[1] wr_data_b[1] ck_en[4] reg_data_4[1] DLH_X1
xi15[0] wr_data_b[0] ck_en[4] reg_data_4[0] DLH_X1
xi7[15] wr_data_b[15] ck_en[0] reg_data_0[15] DLH_X1
xi7[14] wr_data_b[14] ck_en[0] reg_data_0[14] DLH_X1
xi7[13] wr_data_b[13] ck_en[0] reg_data_0[13] DLH_X1
xi7[12] wr_data_b[12] ck_en[0] reg_data_0[12] DLH_X1
xi7[11] wr_data_b[11] ck_en[0] reg_data_0[11] DLH_X1
xi7[10] wr_data_b[10] ck_en[0] reg_data_0[10] DLH_X1
xi7[9] wr_data_b[9] ck_en[0] reg_data_0[9] DLH_X1
xi7[8] wr_data_b[8] ck_en[0] reg_data_0[8] DLH_X1
xi7[7] wr_data_b[7] ck_en[0] reg_data_0[7] DLH_X1
xi7[6] wr_data_b[6] ck_en[0] reg_data_0[6] DLH_X1
xi7[5] wr_data_b[5] ck_en[0] reg_data_0[5] DLH_X1
xi7[4] wr_data_b[4] ck_en[0] reg_data_0[4] DLH_X1
xi7[3] wr_data_b[3] ck_en[0] reg_data_0[3] DLH_X1
xi7[2] wr_data_b[2] ck_en[0] reg_data_0[2] DLH_X1
xi7[1] wr_data_b[1] ck_en[0] reg_data_0[1] DLH_X1
xi7[0] wr_data_b[0] ck_en[0] reg_data_0[0] DLH_X1
xi13[15] wr_data_b[15] ck_en[2] reg_data_2[15] DLH_X1
xi13[14] wr_data_b[14] ck_en[2] reg_data_2[14] DLH_X1
xi13[13] wr_data_b[13] ck_en[2] reg_data_2[13] DLH_X1
xi13[12] wr_data_b[12] ck_en[2] reg_data_2[12] DLH_X1
xi13[11] wr_data_b[11] ck_en[2] reg_data_2[11] DLH_X1
xi13[10] wr_data_b[10] ck_en[2] reg_data_2[10] DLH_X1
xi13[9] wr_data_b[9] ck_en[2] reg_data_2[9] DLH_X1
xi13[8] wr_data_b[8] ck_en[2] reg_data_2[8] DLH_X1
xi13[7] wr_data_b[7] ck_en[2] reg_data_2[7] DLH_X1
xi13[6] wr_data_b[6] ck_en[2] reg_data_2[6] DLH_X1
xi13[5] wr_data_b[5] ck_en[2] reg_data_2[5] DLH_X1
xi13[4] wr_data_b[4] ck_en[2] reg_data_2[4] DLH_X1
xi13[3] wr_data_b[3] ck_en[2] reg_data_2[3] DLH_X1
xi13[2] wr_data_b[2] ck_en[2] reg_data_2[2] DLH_X1
xi13[1] wr_data_b[1] ck_en[2] reg_data_2[1] DLH_X1
xi13[0] wr_data_b[0] ck_en[2] reg_data_2[0] DLH_X1
xi14[15] wr_data_b[15] ck_en[3] reg_data_3[15] DLH_X1
xi14[14] wr_data_b[14] ck_en[3] reg_data_3[14] DLH_X1
xi14[13] wr_data_b[13] ck_en[3] reg_data_3[13] DLH_X1
xi14[12] wr_data_b[12] ck_en[3] reg_data_3[12] DLH_X1
xi14[11] wr_data_b[11] ck_en[3] reg_data_3[11] DLH_X1
xi14[10] wr_data_b[10] ck_en[3] reg_data_3[10] DLH_X1
xi14[9] wr_data_b[9] ck_en[3] reg_data_3[9] DLH_X1
xi14[8] wr_data_b[8] ck_en[3] reg_data_3[8] DLH_X1
xi14[7] wr_data_b[7] ck_en[3] reg_data_3[7] DLH_X1
xi14[6] wr_data_b[6] ck_en[3] reg_data_3[6] DLH_X1
xi14[5] wr_data_b[5] ck_en[3] reg_data_3[5] DLH_X1
xi14[4] wr_data_b[4] ck_en[3] reg_data_3[4] DLH_X1
xi14[3] wr_data_b[3] ck_en[3] reg_data_3[3] DLH_X1
xi14[2] wr_data_b[2] ck_en[3] reg_data_3[2] DLH_X1
xi14[1] wr_data_b[1] ck_en[3] reg_data_3[1] DLH_X1
xi14[0] wr_data_b[0] ck_en[3] reg_data_3[0] DLH_X1
xi8[15] wr_data_b[15] ck_en[1] reg_data_1[15] DLH_X1
xi8[14] wr_data_b[14] ck_en[1] reg_data_1[14] DLH_X1
xi8[13] wr_data_b[13] ck_en[1] reg_data_1[13] DLH_X1
xi8[12] wr_data_b[12] ck_en[1] reg_data_1[12] DLH_X1
xi8[11] wr_data_b[11] ck_en[1] reg_data_1[11] DLH_X1
xi8[10] wr_data_b[10] ck_en[1] reg_data_1[10] DLH_X1
xi8[9] wr_data_b[9] ck_en[1] reg_data_1[9] DLH_X1
xi8[8] wr_data_b[8] ck_en[1] reg_data_1[8] DLH_X1
xi8[7] wr_data_b[7] ck_en[1] reg_data_1[7] DLH_X1
xi8[6] wr_data_b[6] ck_en[1] reg_data_1[6] DLH_X1
xi8[5] wr_data_b[5] ck_en[1] reg_data_1[5] DLH_X1
xi8[4] wr_data_b[4] ck_en[1] reg_data_1[4] DLH_X1
xi8[3] wr_data_b[3] ck_en[1] reg_data_1[3] DLH_X1
xi8[2] wr_data_b[2] ck_en[1] reg_data_1[2] DLH_X1
xi8[1] wr_data_b[1] ck_en[1] reg_data_1[1] DLH_X1
xi8[0] wr_data_b[0] ck_en[1] reg_data_1[0] DLH_X1
.ends cad5_13_16_REGFILE_schematic

.subckt RF 
+ rd_data_0[0] rd_data_0[1] rd_data_0[2] rd_data_0[3] rd_data_0[4] rd_data_0[5] rd_data_0[6] rd_data_0[7]
+ rd_data_0[8] rd_data_0[9] rd_data_0[10] rd_data_0[11] rd_data_0[12] rd_data_0[13] rd_data_0[14] rd_data_0[15]
+ rd_data_1[0] rd_data_1[1] rd_data_1[2] rd_data_1[3] rd_data_1[4] rd_data_1[5] rd_data_1[6] rd_data_1[7]
+ rd_data_1[8] rd_data_1[9] rd_data_1[10] rd_data_1[11] rd_data_1[12] rd_data_1[13] rd_data_1[14] rd_data_1[15]
+ rd_addr_0[0] rd_addr_0[1] rd_addr_0[2] rd_addr_0[3] 
+ rd_addr_1[0] rd_addr_1[1] rd_addr_1[2] rd_addr_1[3] 
+ wr_addr[0] wr_addr[1] wr_addr[2] wr_addr[3] 
+ wr_data[0] wr_data[1] wr_data[2] wr_data[3] wr_data[4] wr_data[5] wr_data[6] wr_data[7]
+ wr_data[8] wr_data[9] wr_data[10] wr_data[11] wr_data[12] wr_data[13] wr_data[14] wr_data[15]
+ wr_en clk
xi1 rd_addr_1[3] rd_addr_1[2] rd_addr_1[1] rd_addr_1[0] r1_d[12] r1_d[11] r1_d[10] r1_d[9] r1_d[8] r1_d[7] r1_d[6] r1_d[5] r1_d[4] r1_d[3] r1_d[2] r1_d[1] r1_d[0] DEC_Read_4_13
xi0 rd_addr_0[3] rd_addr_0[2] rd_addr_0[1] rd_addr_0[0] r0_d[12] r0_d[11] r0_d[10] r0_d[9] r0_d[8] r0_d[7] r0_d[6] r0_d[5] r0_d[4] r0_d[3] r0_d[2] r0_d[1] r0_d[0] DEC_Read_4_13
xi2 clk al_clk_en[12] al_clk_en[11] al_clk_en[10] al_clk_en[9] al_clk_en[8] al_clk_en[7] al_clk_en[6] al_clk_en[5] al_clk_en[4] al_clk_en[3] al_clk_en[2] al_clk_en[1] al_clk_en[0] wr_addr[3] wr_addr[2] wr_addr[1] wr_addr[0] wr_en DEC_EN_4_13
xi3 clk al_clk_en[12] al_clk_en[11] al_clk_en[10] al_clk_en[9] al_clk_en[8] al_clk_en[7] al_clk_en[6] al_clk_en[5] al_clk_en[4] al_clk_en[3] al_clk_en[2] al_clk_en[1] al_clk_en[0] r0_d[12] r0_d[11] r0_d[10] r0_d[9] r0_d[8] r0_d[7] r0_d[6] r0_d[5] r0_d[4] r0_d[3] r0_d[2] r0_d[1] r0_d[0] r1_d[12] r1_d[11] r1_d[10] r1_d[9] r1_d[8] r1_d[7] r1_d[6] r1_d[5] r1_d[4] r1_d[3] r1_d[2] r1_d[1] r1_d[0] rd_data_0[15] rd_data_0[14] rd_data_0[13] rd_data_0[12] rd_data_0[11] rd_data_0[10] rd_data_0[9] rd_data_0[8] rd_data_0[7] rd_data_0[6] rd_data_0[5] rd_data_0[4] rd_data_0[3] rd_data_0[2] rd_data_0[1] rd_data_0[0] rd_data_1[15] rd_data_1[14] rd_data_1[13] rd_data_1[12] rd_data_1[11] rd_data_1[10] rd_data_1[9] rd_data_1[8] rd_data_1[7] rd_data_1[6] rd_data_1[5] rd_data_1[4] rd_data_1[3] rd_data_1[2] rd_data_1[1] rd_data_1[0] wr_data[15] wr_data[14] wr_data[13] wr_data[12] wr_data[11] wr_data[10] wr_data[9] wr_data[8] wr_data[7] wr_data[6] wr_data[5] wr_data[4] wr_data[3] wr_data[2] wr_data[1] wr_data[0] cad5_13_16_REGFILE_schematic
.ends RF
.END
