../part6/ring_osc_2x.ckt