../part4/ring_osc.ckt