** Generated for: hspiceD
** Generated on: Dec  3 16:28:41 2021
** Design library name: cad6
** Design cell name: OUT_MUX_BUF_16B
** Design view name: schematic
.GLOBAL vss! vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad6
** Cell name: MUX2_X1
** View name: schematic
.subckt MUX2_X1 a b s z
m_i_4 net_1 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_5 z_neg x1 net_1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_2 z_neg s net_0 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_3 net_0 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_10 vss! s x1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_6 net_2 s z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_8 vdd! a net_2 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_9 net_3 x1 z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_7 vdd! b net_3 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_11 vdd! s x1 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends MUX2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INV_X1
** View name: schematic
.subckt INV_X1 a zn
m_i_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INV_X4
** View name: schematic
.subckt INV_X4 a zn
m_i_1_0_x4_0 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_1 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_2 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_3 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0_0_x4_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_1 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_2 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_3 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV_X4
** End of subcircuit definition.

** Library name: cad6
** Cell name: BUF_X1
** View name: schematic
.subckt BUF_X1 a z
m_i_3 vdd! a z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_2 vss! a z_neg vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends BUF_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: OUT_MUX_BUF_16B
** View name: schematic
xi0<15> logic_out<15> arithmetic_out<15> ctrl_2_buf<15> alu_pre<15> MUX2_X1
xi0<14> logic_out<14> arithmetic_out<14> ctrl_2_buf<14> alu_pre<14> MUX2_X1
xi0<13> logic_out<13> arithmetic_out<13> ctrl_2_buf<13> alu_pre<13> MUX2_X1
xi0<12> logic_out<12> arithmetic_out<12> ctrl_2_buf<12> alu_pre<12> MUX2_X1
xi0<11> logic_out<11> arithmetic_out<11> ctrl_2_buf<11> alu_pre<11> MUX2_X1
xi0<10> logic_out<10> arithmetic_out<10> ctrl_2_buf<10> alu_pre<10> MUX2_X1
xi0<9> logic_out<9> arithmetic_out<9> ctrl_2_buf<9> alu_pre<9> MUX2_X1
xi0<8> logic_out<8> arithmetic_out<8> ctrl_2_buf<8> alu_pre<8> MUX2_X1
xi0<7> logic_out<7> arithmetic_out<7> ctrl_2_buf<7> alu_pre<7> MUX2_X1
xi0<6> logic_out<6> arithmetic_out<6> ctrl_2_buf<6> alu_pre<6> MUX2_X1
xi0<5> logic_out<5> arithmetic_out<5> ctrl_2_buf<5> alu_pre<5> MUX2_X1
xi0<4> logic_out<4> arithmetic_out<4> ctrl_2_buf<4> alu_pre<4> MUX2_X1
xi0<3> logic_out<3> arithmetic_out<3> ctrl_2_buf<3> alu_pre<3> MUX2_X1
xi0<2> logic_out<2> arithmetic_out<2> ctrl_2_buf<2> alu_pre<2> MUX2_X1
xi0<1> logic_out<1> arithmetic_out<1> ctrl_2_buf<1> alu_pre<1> MUX2_X1
xi0<0> logic_out<0> arithmetic_out<0> ctrl_2_buf<0> alu_pre<0> MUX2_X1
xi1<15> alu_pre<15> net3<0> INV_X1
xi1<14> alu_pre<14> net3<1> INV_X1
xi1<13> alu_pre<13> net3<2> INV_X1
xi1<12> alu_pre<12> net3<3> INV_X1
xi1<11> alu_pre<11> net3<4> INV_X1
xi1<10> alu_pre<10> net3<5> INV_X1
xi1<9> alu_pre<9> net3<6> INV_X1
xi1<8> alu_pre<8> net3<7> INV_X1
xi1<7> alu_pre<7> net3<8> INV_X1
xi1<6> alu_pre<6> net3<9> INV_X1
xi1<5> alu_pre<5> net3<10> INV_X1
xi1<4> alu_pre<4> net3<11> INV_X1
xi1<3> alu_pre<3> net3<12> INV_X1
xi1<2> alu_pre<2> net3<13> INV_X1
xi1<1> alu_pre<1> net3<14> INV_X1
xi1<0> alu_pre<0> net3<15> INV_X1
xi2<15> net3<0> alu_out<15> INV_X4
xi2<14> net3<1> alu_out<14> INV_X4
xi2<13> net3<2> alu_out<13> INV_X4
xi2<12> net3<3> alu_out<12> INV_X4
xi2<11> net3<4> alu_out<11> INV_X4
xi2<10> net3<5> alu_out<10> INV_X4
xi2<9> net3<6> alu_out<9> INV_X4
xi2<8> net3<7> alu_out<8> INV_X4
xi2<7> net3<8> alu_out<7> INV_X4
xi2<6> net3<9> alu_out<6> INV_X4
xi2<5> net3<10> alu_out<5> INV_X4
xi2<4> net3<11> alu_out<4> INV_X4
xi2<3> net3<12> alu_out<3> INV_X4
xi2<2> net3<13> alu_out<2> INV_X4
xi2<1> net3<14> alu_out<1> INV_X4
xi2<0> net3<15> alu_out<0> INV_X4
xi27 ctrl_2_buf<13> ctrl_2_buf<12> BUF_X1
xi26 ctrl_2_buf<14> ctrl_2_buf<13> BUF_X1
xi25 ctrl_2_buf<15> ctrl_2_buf<14> BUF_X1
xi24 ctrl<2> ctrl_2_buf<15> BUF_X1
xi23 ctrl_2_buf<12> ctrl_2_buf<11> BUF_X1
xi22 ctrl_2_buf<11> ctrl_2_buf<10> BUF_X1
xi21 ctrl_2_buf<10> ctrl_2_buf<9> BUF_X1
xi20 ctrl_2_buf<9> ctrl_2_buf<8> BUF_X1
xi19 ctrl_2_buf<5> ctrl_2_buf<4> BUF_X1
xi18 ctrl_2_buf<6> ctrl_2_buf<5> BUF_X1
xi17 ctrl_2_buf<7> ctrl_2_buf<6> BUF_X1
xi16 ctrl_2_buf<8> ctrl_2_buf<7> BUF_X1
xi12 ctrl_2_buf<4> ctrl_2_buf<3> BUF_X1
xi11 ctrl_2_buf<3> ctrl_2_buf<2> BUF_X1
xi4 ctrl_2_buf<2> ctrl_2_buf<1> BUF_X1
xi3 ctrl_2_buf<1> ctrl_2_buf<0> BUF_X1
.END
