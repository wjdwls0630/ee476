.GLOBAL vss! vdd!


.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2

.subckt NAND2_balanced a b z W=500e-9
mnmos1 net2 b vss! vss! NMOS_VTG L=60e-9 W=350e-9 AD=36.75e-15 AS=36.75e-15 PD=560e-9 PS=560e-9 M=1
mnmos0 z a net2 vss! NMOS_VTG L=60e-9 W=350e-9 AD=36.75e-15 AS=36.75e-15 PD=560e-9 PS=560e-9 M=1
mpmos1 z b vdd! vdd! PMOS_VTG L=60e-9 W='W' AD='0.105e-6*W' AS='0.105e-6*W' PD='W+210e-9' PS='W+210e-9' M=1
mpmos0 z a vdd! vdd! PMOS_VTG L=60e-9 W='W' AD='0.105e-6*W' AS='0.105e-6*W' PD='W+210e-9' PS='W+210e-9' M=1
.ends NAND2_balanced

