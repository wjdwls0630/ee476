* File: RF.pex.netlist
* Created: Mon Nov 22 22:20:54 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.GLOBAL vdd! vss!

.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

.subckt RF 
+ rd_data_0<0> rd_data_0<1> rd_data_0<2> rd_data_0<3> rd_data_0<4> rd_data_0<5> rd_data_0<6> rd_data_0<7>
+ rd_data_0<8> rd_data_0<9> rd_data_0<10> rd_data_0<11> rd_data_0<12> rd_data_0<13> rd_data_0<14> rd_data_0<15>
+ rd_data_1<0> rd_data_1<1> rd_data_1<2> rd_data_1<3> rd_data_1<4> rd_data_1<5> rd_data_1<6> rd_data_1<7>
+ rd_data_1<8> rd_data_1<9> rd_data_1<10> rd_data_1<11> rd_data_1<12> rd_data_1<13> rd_data_1<14> rd_data_1<15>
+ rd_addr_0<0> rd_addr_0<1> rd_addr_0<2> rd_addr_0<3> 
+ rd_addr_1<0> rd_addr_1<1> rd_addr_1<2> rd_addr_1<3> 
+ wr_addr<0> wr_addr<1> wr_addr<2> wr_addr<3> 
+ wr_data<0> wr_data<1> wr_data<2> wr_data<3> wr_data<4> wr_data<5> wr_data<6> wr_data<7>
+ wr_data<8> wr_data<9> wr_data<10> wr_data<11> wr_data<12> wr_data<13> wr_data<14> wr_data<15>
+ wr_en clk
* 
mXI0.XI0.XI24.MM_i_1 XI0.XI0.XI24.NET_0 XI0.XI0.NET_11XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI24.MM_i_0 XI0.NET1<0> XI0.XI0.NET_XX00 XI0.XI0.XI24.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI24.MM_i_3 XI0.NET1<0> XI0.XI0.NET_11XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI24.MM_i_2 VDD! XI0.XI0.NET_XX00 XI0.NET1<0> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI23.MM_i_1 XI0.XI0.XI23.NET_0 XI0.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI23.MM_i_0 XI0.NET1<1> XI0.XI0.NET_XX11 XI0.XI0.XI23.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI23.MM_i_3 XI0.NET1<1> XI0.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI23.MM_i_2 VDD! XI0.XI0.NET_XX11 XI0.NET1<1> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI22.MM_i_1 XI0.XI0.XI22.NET_0 XI0.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI22.MM_i_0 XI0.NET1<2> XI0.XI0.NET_XX10 XI0.XI0.XI22.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI22.MM_i_3 XI0.NET1<2> XI0.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI22.MM_i_2 VDD! XI0.XI0.NET_XX10 XI0.NET1<2> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI21.MM_i_1 XI0.XI0.XI21.NET_0 XI0.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI21.MM_i_0 XI0.NET1<3> XI0.XI0.NET_XX01 XI0.XI0.XI21.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI21.MM_i_3 XI0.NET1<3> XI0.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI21.MM_i_2 VDD! XI0.XI0.NET_XX01 XI0.NET1<3> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI20.MM_i_1 XI0.XI0.XI20.NET_0 XI0.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI20.MM_i_0 XI0.NET1<4> XI0.XI0.NET_XX00 XI0.XI0.XI20.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI20.MM_i_3 XI0.NET1<4> XI0.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI20.MM_i_2 VDD! XI0.XI0.NET_XX00 XI0.NET1<4> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI19.MM_i_1 XI0.XI0.XI19.NET_0 XI0.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI19.MM_i_0 XI0.NET1<5> XI0.XI0.NET_XX11 XI0.XI0.XI19.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI19.MM_i_3 XI0.NET1<5> XI0.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI19.MM_i_2 VDD! XI0.XI0.NET_XX11 XI0.NET1<5> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI18.MM_i_1 XI0.XI0.XI18.NET_0 XI0.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI18.MM_i_0 XI0.NET1<6> XI0.XI0.NET_XX10 XI0.XI0.XI18.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI18.MM_i_3 XI0.NET1<6> XI0.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI18.MM_i_2 VDD! XI0.XI0.NET_XX10 XI0.NET1<6> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI17.MM_i_1 XI0.XI0.XI17.NET_0 XI0.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI17.MM_i_0 XI0.NET1<7> XI0.XI0.NET_XX01 XI0.XI0.XI17.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI17.MM_i_3 XI0.NET1<7> XI0.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI17.MM_i_2 VDD! XI0.XI0.NET_XX01 XI0.NET1<7> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI16.MM_i_1 XI0.XI0.XI16.NET_0 XI0.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI16.MM_i_0 XI0.NET1<8> XI0.XI0.NET_XX00 XI0.XI0.XI16.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI16.MM_i_3 XI0.NET1<8> XI0.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI16.MM_i_2 VDD! XI0.XI0.NET_XX00 XI0.NET1<8> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI15.MM_i_1 XI0.XI0.XI15.NET_0 XI0.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI15.MM_i_0 XI0.NET1<9> XI0.XI0.NET_XX11 XI0.XI0.XI15.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI15.MM_i_3 XI0.NET1<9> XI0.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI15.MM_i_2 VDD! XI0.XI0.NET_XX11 XI0.NET1<9> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI14.MM_i_1 XI0.XI0.XI14.NET_0 XI0.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI14.MM_i_0 XI0.NET1<10> XI0.XI0.NET_XX10 XI0.XI0.XI14.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI14.MM_i_3 XI0.NET1<10> XI0.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI14.MM_i_2 VDD! XI0.XI0.NET_XX10 XI0.NET1<10> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI13.MM_i_1 XI0.XI0.XI13.NET_0 XI0.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI13.MM_i_0 XI0.NET1<11> XI0.XI0.NET_XX01 XI0.XI0.XI13.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI13.MM_i_3 XI0.NET1<11> XI0.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI13.MM_i_2 VDD! XI0.XI0.NET_XX01 XI0.NET1<11> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI12.MM_i_1 XI0.XI0.XI12.NET_0 XI0.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI0.XI12.MM_i_0 XI0.NET1<12> XI0.XI0.NET_XX00 XI0.XI0.XI12.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI12.MM_i_3 XI0.NET1<12> XI0.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI0.XI12.MM_i_2 VDD! XI0.XI0.NET_XX00 XI0.NET1<12> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI11.MM_i_2 XI0.XI0.XI11.NET_0 RD_ADDR_0<2> XI0.XI0.XI11.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI11.MM_i_3 VSS! RD_ADDR_0<3> XI0.XI0.XI11.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI11.MM_i_0 XI0.XI0.NET_11XX XI0.XI0.XI11.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI11.MM_i_4 XI0.XI0.XI11.ZN_NEG RD_ADDR_0<2> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI11.MM_i_5 VDD! RD_ADDR_0<3> XI0.XI0.XI11.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI11.MM_i_1 XI0.XI0.NET_11XX XI0.XI0.XI11.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI7.MM_i_2 XI0.XI0.XI7.NET_0 RD_ADDR_0<0> XI0.XI0.XI7.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI7.MM_i_3 VSS! RD_ADDR_0<1> XI0.XI0.XI7.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI7.MM_i_0 XI0.XI0.NET_XX11 XI0.XI0.XI7.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI7.MM_i_4 XI0.XI0.XI7.ZN_NEG RD_ADDR_0<0> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI7.MM_i_5 VDD! RD_ADDR_0<1> XI0.XI0.XI7.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI7.MM_i_1 XI0.XI0.NET_XX11 XI0.XI0.XI7.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI10.MM_i_2 XI0.XI0.XI10.NET_0 XI0.XI0.ADDR_BAR<2> XI0.XI0.XI10.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI10.MM_i_3 VSS! RD_ADDR_0<3> XI0.XI0.XI10.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI10.MM_i_0 XI0.XI0.NET_10XX XI0.XI0.XI10.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI10.MM_i_4 XI0.XI0.XI10.ZN_NEG XI0.XI0.ADDR_BAR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI10.MM_i_5 VDD! RD_ADDR_0<3> XI0.XI0.XI10.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI10.MM_i_1 XI0.XI0.NET_10XX XI0.XI0.XI10.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI6.MM_i_2 XI0.XI0.XI6.NET_0 XI0.XI0.ADDR_BAR<0> XI0.XI0.XI6.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI6.MM_i_3 VSS! RD_ADDR_0<1> XI0.XI0.XI6.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI6.MM_i_0 XI0.XI0.NET_XX10 XI0.XI0.XI6.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI6.MM_i_4 XI0.XI0.XI6.ZN_NEG XI0.XI0.ADDR_BAR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI6.MM_i_5 VDD! RD_ADDR_0<1> XI0.XI0.XI6.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI6.MM_i_1 XI0.XI0.NET_XX10 XI0.XI0.XI6.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI9.MM_i_2 XI0.XI0.XI9.NET_0 RD_ADDR_0<2> XI0.XI0.XI9.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI9.MM_i_3 VSS! XI0.XI0.ADDR_BAR<3> XI0.XI0.XI9.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI9.MM_i_0 XI0.XI0.NET_01XX XI0.XI0.XI9.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI9.MM_i_4 XI0.XI0.XI9.ZN_NEG RD_ADDR_0<2> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI9.MM_i_5 VDD! XI0.XI0.ADDR_BAR<3> XI0.XI0.XI9.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI9.MM_i_1 XI0.XI0.NET_01XX XI0.XI0.XI9.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI5.MM_i_2 XI0.XI0.XI5.NET_0 RD_ADDR_0<0> XI0.XI0.XI5.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI5.MM_i_3 VSS! XI0.XI0.ADDR_BAR<1> XI0.XI0.XI5.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI5.MM_i_0 XI0.XI0.NET_XX01 XI0.XI0.XI5.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI5.MM_i_4 XI0.XI0.XI5.ZN_NEG RD_ADDR_0<0> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI5.MM_i_5 VDD! XI0.XI0.ADDR_BAR<1> XI0.XI0.XI5.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI5.MM_i_1 XI0.XI0.NET_XX01 XI0.XI0.XI5.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI8.MM_i_2 XI0.XI0.XI8.NET_0 XI0.XI0.ADDR_BAR<2> XI0.XI0.XI8.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI8.MM_i_3 VSS! XI0.XI0.ADDR_BAR<3> XI0.XI0.XI8.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI8.MM_i_0 XI0.XI0.NET_00XX XI0.XI0.XI8.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI8.MM_i_4 XI0.XI0.XI8.ZN_NEG XI0.XI0.ADDR_BAR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI8.MM_i_5 VDD! XI0.XI0.ADDR_BAR<3> XI0.XI0.XI8.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI8.MM_i_1 XI0.XI0.NET_00XX XI0.XI0.XI8.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI4.MM_i_2 XI0.XI0.XI4.NET_0 XI0.XI0.ADDR_BAR<0> XI0.XI0.XI4.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI0.XI0.XI4.MM_i_3 VSS! XI0.XI0.ADDR_BAR<1> XI0.XI0.XI4.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI0.XI0.XI4.MM_i_0 XI0.XI0.NET_XX00 XI0.XI0.XI4.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI0.XI4.MM_i_4 XI0.XI0.XI4.ZN_NEG XI0.XI0.ADDR_BAR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI0.XI0.XI4.MM_i_5 VDD! XI0.XI0.ADDR_BAR<1> XI0.XI0.XI4.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI0.XI0.XI4.MM_i_1 XI0.XI0.NET_XX00 XI0.XI0.XI4.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI0.XI0.XI2.MM_i_0 XI0.XI0.ADDR_BAR<2> RD_ADDR_0<2> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI0.XI0.XI2.MM_i_1 XI0.XI0.ADDR_BAR<2> RD_ADDR_0<2> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI0.XI0.XI0.MM_i_0 XI0.XI0.ADDR_BAR<0> RD_ADDR_0<0> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI0.XI0.XI0.MM_i_1 XI0.XI0.ADDR_BAR<0> RD_ADDR_0<0> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI0.XI0.XI3.MM_i_0 XI0.XI0.ADDR_BAR<3> RD_ADDR_0<3> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI0.XI0.XI3.MM_i_1 XI0.XI0.ADDR_BAR<3> RD_ADDR_0<3> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI0.XI0.XI1.MM_i_0 XI0.XI0.ADDR_BAR<1> RD_ADDR_0<1> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI0.XI0.XI1.MM_i_1 XI0.XI0.ADDR_BAR<1> RD_ADDR_0<1> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<3>.MM_i_0 VSS! XI0.XI1.XI15.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<3>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<3>.MM_i_0_15 VSS! REG_DATA_0<3> XI0.XI1.XI15.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<3>.MM_i_0_15_63 XI0.XI1.XI15.XI3<3>.DUMMY1 REG_DATA_0<3>
+ XI0.XI1.XI15.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<3>.NEN
+ XI0.XI1.XI15.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<3>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<3>.MM_i_24 VDD! XI0.XI1.XI15.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<3>.MM_i_24_1 XI0.XI1.XI15.XI3<3>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<3>.MM_i_24_0 VDD! REG_DATA_0<3> XI0.XI1.XI15.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_0<3> XI0.XI1.XI15.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<3>.MM_i_24_1_48 XI0.XI1.XI15.XI3<3>.Y XI0.XI1.XI15.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<3>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<2>.MM_i_0 VSS! XI0.XI1.XI15.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<2>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<2>.MM_i_0_15 VSS! REG_DATA_0<2> XI0.XI1.XI15.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<2>.MM_i_0_15_63 XI0.XI1.XI15.XI3<2>.DUMMY1 REG_DATA_0<2>
+ XI0.XI1.XI15.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<2>.NEN
+ XI0.XI1.XI15.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<2>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<2>.MM_i_24 VDD! XI0.XI1.XI15.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<2>.MM_i_24_1 XI0.XI1.XI15.XI3<2>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<2>.MM_i_24_0 VDD! REG_DATA_0<2> XI0.XI1.XI15.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_0<2> XI0.XI1.XI15.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<2>.MM_i_24_1_48 XI0.XI1.XI15.XI3<2>.Y XI0.XI1.XI15.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<2>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<1>.MM_i_0 VSS! XI0.XI1.XI15.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<1>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<1>.MM_i_0_15 VSS! REG_DATA_0<1> XI0.XI1.XI15.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<1>.MM_i_0_15_63 XI0.XI1.XI15.XI3<1>.DUMMY1 REG_DATA_0<1>
+ XI0.XI1.XI15.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<1>.NEN
+ XI0.XI1.XI15.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<1>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<1>.MM_i_24 VDD! XI0.XI1.XI15.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<1>.MM_i_24_1 XI0.XI1.XI15.XI3<1>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<1>.MM_i_24_0 VDD! REG_DATA_0<1> XI0.XI1.XI15.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_0<1> XI0.XI1.XI15.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<1>.MM_i_24_1_48 XI0.XI1.XI15.XI3<1>.Y XI0.XI1.XI15.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<1>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<0>.MM_i_0 VSS! XI0.XI1.XI15.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<0>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<0>.MM_i_0_15 VSS! REG_DATA_0<0> XI0.XI1.XI15.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<0>.MM_i_0_15_63 XI0.XI1.XI15.XI3<0>.DUMMY1 REG_DATA_0<0>
+ XI0.XI1.XI15.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<0>.NEN
+ XI0.XI1.XI15.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<0>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<0>.MM_i_24 VDD! XI0.XI1.XI15.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<0>.MM_i_24_1 XI0.XI1.XI15.XI3<0>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<0>.MM_i_24_0 VDD! REG_DATA_0<0> XI0.XI1.XI15.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_0<0> XI0.XI1.XI15.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<0>.MM_i_24_1_48 XI0.XI1.XI15.XI3<0>.Y XI0.XI1.XI15.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<0>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<7>.MM_i_0 VSS! XI0.XI1.XI15.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<7>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<7>.MM_i_0_15 VSS! REG_DATA_0<7> XI0.XI1.XI15.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<7>.MM_i_0_15_63 XI0.XI1.XI15.XI3<7>.DUMMY1 REG_DATA_0<7>
+ XI0.XI1.XI15.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<7>.NEN
+ XI0.XI1.XI15.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<7>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<7>.MM_i_24 VDD! XI0.XI1.XI15.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<7>.MM_i_24_1 XI0.XI1.XI15.XI3<7>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<7>.MM_i_24_0 VDD! REG_DATA_0<7> XI0.XI1.XI15.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_0<7> XI0.XI1.XI15.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<7>.MM_i_24_1_48 XI0.XI1.XI15.XI3<7>.Y XI0.XI1.XI15.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<7>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<6>.MM_i_0 VSS! XI0.XI1.XI15.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<6>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<6>.MM_i_0_15 VSS! REG_DATA_0<6> XI0.XI1.XI15.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<6>.MM_i_0_15_63 XI0.XI1.XI15.XI3<6>.DUMMY1 REG_DATA_0<6>
+ XI0.XI1.XI15.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<6>.NEN
+ XI0.XI1.XI15.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<6>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<6>.MM_i_24 VDD! XI0.XI1.XI15.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<6>.MM_i_24_1 XI0.XI1.XI15.XI3<6>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<6>.MM_i_24_0 VDD! REG_DATA_0<6> XI0.XI1.XI15.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_0<6> XI0.XI1.XI15.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<6>.MM_i_24_1_48 XI0.XI1.XI15.XI3<6>.Y XI0.XI1.XI15.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<6>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<5>.MM_i_0 VSS! XI0.XI1.XI15.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<5>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<5>.MM_i_0_15 VSS! REG_DATA_0<5> XI0.XI1.XI15.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<5>.MM_i_0_15_63 XI0.XI1.XI15.XI3<5>.DUMMY1 REG_DATA_0<5>
+ XI0.XI1.XI15.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<5>.NEN
+ XI0.XI1.XI15.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<5>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<5>.MM_i_24 VDD! XI0.XI1.XI15.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<5>.MM_i_24_1 XI0.XI1.XI15.XI3<5>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<5>.MM_i_24_0 VDD! REG_DATA_0<5> XI0.XI1.XI15.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_0<5> XI0.XI1.XI15.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<5>.MM_i_24_1_48 XI0.XI1.XI15.XI3<5>.Y XI0.XI1.XI15.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<5>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<4>.MM_i_0 VSS! XI0.XI1.XI15.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<4>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<4>.MM_i_0_15 VSS! REG_DATA_0<4> XI0.XI1.XI15.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<4>.MM_i_0_15_63 XI0.XI1.XI15.XI3<4>.DUMMY1 REG_DATA_0<4>
+ XI0.XI1.XI15.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<4>.NEN
+ XI0.XI1.XI15.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<4>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<4>.MM_i_24 VDD! XI0.XI1.XI15.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<4>.MM_i_24_1 XI0.XI1.XI15.XI3<4>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<4>.MM_i_24_0 VDD! REG_DATA_0<4> XI0.XI1.XI15.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_0<4> XI0.XI1.XI15.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<4>.MM_i_24_1_48 XI0.XI1.XI15.XI3<4>.Y XI0.XI1.XI15.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<4>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<11>.MM_i_0 VSS! XI0.XI1.XI15.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<11>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<11>.MM_i_0_15 VSS! REG_DATA_0<11> XI0.XI1.XI15.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<11>.MM_i_0_15_63 XI0.XI1.XI15.XI3<11>.DUMMY1 REG_DATA_0<11>
+ XI0.XI1.XI15.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<11>.NEN
+ XI0.XI1.XI15.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<11>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<11>.MM_i_24 VDD! XI0.XI1.XI15.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<11>.MM_i_24_1 XI0.XI1.XI15.XI3<11>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<11>.MM_i_24_0 VDD! REG_DATA_0<11> XI0.XI1.XI15.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_0<11> XI0.XI1.XI15.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<11>.MM_i_24_1_48 XI0.XI1.XI15.XI3<11>.Y
+ XI0.XI1.XI15.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI15.XI3<11>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<10>.MM_i_0 VSS! XI0.XI1.XI15.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<10>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<10>.MM_i_0_15 VSS! REG_DATA_0<10> XI0.XI1.XI15.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<10>.MM_i_0_15_63 XI0.XI1.XI15.XI3<10>.DUMMY1 REG_DATA_0<10>
+ XI0.XI1.XI15.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<10>.NEN
+ XI0.XI1.XI15.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<10>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<10>.MM_i_24 VDD! XI0.XI1.XI15.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<10>.MM_i_24_1 XI0.XI1.XI15.XI3<10>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<10>.MM_i_24_0 VDD! REG_DATA_0<10> XI0.XI1.XI15.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_0<10> XI0.XI1.XI15.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<10>.MM_i_24_1_48 XI0.XI1.XI15.XI3<10>.Y
+ XI0.XI1.XI15.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI15.XI3<10>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<9>.MM_i_0 VSS! XI0.XI1.XI15.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<9>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<9>.MM_i_0_15 VSS! REG_DATA_0<9> XI0.XI1.XI15.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<9>.MM_i_0_15_63 XI0.XI1.XI15.XI3<9>.DUMMY1 REG_DATA_0<9>
+ XI0.XI1.XI15.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<9>.NEN
+ XI0.XI1.XI15.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<9>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<9>.MM_i_24 VDD! XI0.XI1.XI15.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<9>.MM_i_24_1 XI0.XI1.XI15.XI3<9>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<9>.MM_i_24_0 VDD! REG_DATA_0<9> XI0.XI1.XI15.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_0<9> XI0.XI1.XI15.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<9>.MM_i_24_1_48 XI0.XI1.XI15.XI3<9>.Y XI0.XI1.XI15.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<9>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<8>.MM_i_0 VSS! XI0.XI1.XI15.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<8>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<8>.MM_i_0_15 VSS! REG_DATA_0<8> XI0.XI1.XI15.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<8>.MM_i_0_15_63 XI0.XI1.XI15.XI3<8>.DUMMY1 REG_DATA_0<8>
+ XI0.XI1.XI15.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<8>.NEN
+ XI0.XI1.XI15.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<8>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<8>.MM_i_24 VDD! XI0.XI1.XI15.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<8>.MM_i_24_1 XI0.XI1.XI15.XI3<8>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<8>.MM_i_24_0 VDD! REG_DATA_0<8> XI0.XI1.XI15.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_0<8> XI0.XI1.XI15.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI15.XI3<8>.MM_i_24_1_48 XI0.XI1.XI15.XI3<8>.Y XI0.XI1.XI15.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI15.XI3<8>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<15>.MM_i_0 VSS! XI0.XI1.XI15.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<15>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<15>.MM_i_0_15 VSS! REG_DATA_0<15> XI0.XI1.XI15.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<15>.MM_i_0_15_63 XI0.XI1.XI15.XI3<15>.DUMMY1 REG_DATA_0<15>
+ XI0.XI1.XI15.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<15>.NEN
+ XI0.XI1.XI15.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<15>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<15>.MM_i_24 VDD! XI0.XI1.XI15.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<15>.MM_i_24_1 XI0.XI1.XI15.XI3<15>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<15>.MM_i_24_0 VDD! REG_DATA_0<15> XI0.XI1.XI15.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_0<15> XI0.XI1.XI15.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<15>.MM_i_24_1_48 XI0.XI1.XI15.XI3<15>.Y
+ XI0.XI1.XI15.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI15.XI3<15>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<14>.MM_i_0 VSS! XI0.XI1.XI15.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<14>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<14>.MM_i_0_15 VSS! REG_DATA_0<14> XI0.XI1.XI15.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<14>.MM_i_0_15_63 XI0.XI1.XI15.XI3<14>.DUMMY1 REG_DATA_0<14>
+ XI0.XI1.XI15.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<14>.NEN
+ XI0.XI1.XI15.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<14>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<14>.MM_i_24 VDD! XI0.XI1.XI15.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<14>.MM_i_24_1 XI0.XI1.XI15.XI3<14>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<14>.MM_i_24_0 VDD! REG_DATA_0<14> XI0.XI1.XI15.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_0<14> XI0.XI1.XI15.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<14>.MM_i_24_1_48 XI0.XI1.XI15.XI3<14>.Y
+ XI0.XI1.XI15.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI15.XI3<14>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<13>.MM_i_0 VSS! XI0.XI1.XI15.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<13>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<13>.MM_i_0_15 VSS! REG_DATA_0<13> XI0.XI1.XI15.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<13>.MM_i_0_15_63 XI0.XI1.XI15.XI3<13>.DUMMY1 REG_DATA_0<13>
+ XI0.XI1.XI15.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<13>.NEN
+ XI0.XI1.XI15.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<13>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<13>.MM_i_24 VDD! XI0.XI1.XI15.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<13>.MM_i_24_1 XI0.XI1.XI15.XI3<13>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<13>.MM_i_24_0 VDD! REG_DATA_0<13> XI0.XI1.XI15.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_0<13> XI0.XI1.XI15.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<13>.MM_i_24_1_48 XI0.XI1.XI15.XI3<13>.Y
+ XI0.XI1.XI15.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI15.XI3<13>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI15.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI15.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI15.XI3<12>.MM_i_0 VSS! XI0.XI1.XI15.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI15.XI3<12>.MM_i_0_14 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<12>.MM_i_0_15 VSS! REG_DATA_0<12> XI0.XI1.XI15.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<12>.MM_i_0_15_63 XI0.XI1.XI15.XI3<12>.DUMMY1 REG_DATA_0<12>
+ XI0.XI1.XI15.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI15.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI15.XI3<12>.NEN
+ XI0.XI1.XI15.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI15.XI3<12>.MM_i_17 VSS! XI0.NET1<12> XI0.XI1.XI15.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI15.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI15.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<12>.MM_i_24 VDD! XI0.XI1.XI15.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI15.XI3<12>.MM_i_24_1 XI0.XI1.XI15.XI3<12>.DUMMY0 XI0.NET1<12>
+ XI0.XI1.XI15.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI15.XI3<12>.MM_i_24_0 VDD! REG_DATA_0<12> XI0.XI1.XI15.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_0<12> XI0.XI1.XI15.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI15.XI3<12>.MM_i_24_1_48 XI0.XI1.XI15.XI3<12>.Y
+ XI0.XI1.XI15.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI15.XI3<12>.MM_i_42 VDD! XI0.NET1<12> XI0.XI1.XI15.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<3>.MM_i_0 VSS! XI0.XI1.XI3.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<3>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<3>.MM_i_0_15 VSS! REG_DATA_12<3> XI0.XI1.XI3.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<3>.MM_i_0_15_63 XI0.XI1.XI3.XI3<3>.DUMMY1 REG_DATA_12<3>
+ XI0.XI1.XI3.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<3>.NEN
+ XI0.XI1.XI3.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<3>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<3>.MM_i_24 VDD! XI0.XI1.XI3.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<3>.MM_i_24_1 XI0.XI1.XI3.XI3<3>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<3>.MM_i_24_0 VDD! REG_DATA_12<3> XI0.XI1.XI3.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_12<3> XI0.XI1.XI3.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<3>.MM_i_24_1_48 XI0.XI1.XI3.XI3<3>.Y XI0.XI1.XI3.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<3>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<2>.MM_i_0 VSS! XI0.XI1.XI3.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<2>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<2>.MM_i_0_15 VSS! REG_DATA_12<2> XI0.XI1.XI3.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<2>.MM_i_0_15_63 XI0.XI1.XI3.XI3<2>.DUMMY1 REG_DATA_12<2>
+ XI0.XI1.XI3.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<2>.NEN
+ XI0.XI1.XI3.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<2>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<2>.MM_i_24 VDD! XI0.XI1.XI3.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<2>.MM_i_24_1 XI0.XI1.XI3.XI3<2>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<2>.MM_i_24_0 VDD! REG_DATA_12<2> XI0.XI1.XI3.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_12<2> XI0.XI1.XI3.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<2>.MM_i_24_1_48 XI0.XI1.XI3.XI3<2>.Y XI0.XI1.XI3.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<2>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<1>.MM_i_0 VSS! XI0.XI1.XI3.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<1>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<1>.MM_i_0_15 VSS! REG_DATA_12<1> XI0.XI1.XI3.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<1>.MM_i_0_15_63 XI0.XI1.XI3.XI3<1>.DUMMY1 REG_DATA_12<1>
+ XI0.XI1.XI3.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<1>.NEN
+ XI0.XI1.XI3.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<1>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<1>.MM_i_24 VDD! XI0.XI1.XI3.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<1>.MM_i_24_1 XI0.XI1.XI3.XI3<1>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<1>.MM_i_24_0 VDD! REG_DATA_12<1> XI0.XI1.XI3.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_12<1> XI0.XI1.XI3.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<1>.MM_i_24_1_48 XI0.XI1.XI3.XI3<1>.Y XI0.XI1.XI3.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<1>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<0>.MM_i_0 VSS! XI0.XI1.XI3.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<0>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<0>.MM_i_0_15 VSS! REG_DATA_12<0> XI0.XI1.XI3.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<0>.MM_i_0_15_63 XI0.XI1.XI3.XI3<0>.DUMMY1 REG_DATA_12<0>
+ XI0.XI1.XI3.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<0>.NEN
+ XI0.XI1.XI3.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<0>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<0>.MM_i_24 VDD! XI0.XI1.XI3.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<0>.MM_i_24_1 XI0.XI1.XI3.XI3<0>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<0>.MM_i_24_0 VDD! REG_DATA_12<0> XI0.XI1.XI3.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_12<0> XI0.XI1.XI3.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<0>.MM_i_24_1_48 XI0.XI1.XI3.XI3<0>.Y XI0.XI1.XI3.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<0>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<7>.MM_i_0 VSS! XI0.XI1.XI3.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<7>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<7>.MM_i_0_15 VSS! REG_DATA_12<7> XI0.XI1.XI3.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<7>.MM_i_0_15_63 XI0.XI1.XI3.XI3<7>.DUMMY1 REG_DATA_12<7>
+ XI0.XI1.XI3.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<7>.NEN
+ XI0.XI1.XI3.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<7>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<7>.MM_i_24 VDD! XI0.XI1.XI3.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<7>.MM_i_24_1 XI0.XI1.XI3.XI3<7>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<7>.MM_i_24_0 VDD! REG_DATA_12<7> XI0.XI1.XI3.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_12<7> XI0.XI1.XI3.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<7>.MM_i_24_1_48 XI0.XI1.XI3.XI3<7>.Y XI0.XI1.XI3.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<7>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<6>.MM_i_0 VSS! XI0.XI1.XI3.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<6>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<6>.MM_i_0_15 VSS! REG_DATA_12<6> XI0.XI1.XI3.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<6>.MM_i_0_15_63 XI0.XI1.XI3.XI3<6>.DUMMY1 REG_DATA_12<6>
+ XI0.XI1.XI3.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<6>.NEN
+ XI0.XI1.XI3.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<6>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<6>.MM_i_24 VDD! XI0.XI1.XI3.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<6>.MM_i_24_1 XI0.XI1.XI3.XI3<6>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<6>.MM_i_24_0 VDD! REG_DATA_12<6> XI0.XI1.XI3.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_12<6> XI0.XI1.XI3.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<6>.MM_i_24_1_48 XI0.XI1.XI3.XI3<6>.Y XI0.XI1.XI3.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<6>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<5>.MM_i_0 VSS! XI0.XI1.XI3.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<5>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<5>.MM_i_0_15 VSS! REG_DATA_12<5> XI0.XI1.XI3.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<5>.MM_i_0_15_63 XI0.XI1.XI3.XI3<5>.DUMMY1 REG_DATA_12<5>
+ XI0.XI1.XI3.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<5>.NEN
+ XI0.XI1.XI3.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<5>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<5>.MM_i_24 VDD! XI0.XI1.XI3.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<5>.MM_i_24_1 XI0.XI1.XI3.XI3<5>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<5>.MM_i_24_0 VDD! REG_DATA_12<5> XI0.XI1.XI3.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_12<5> XI0.XI1.XI3.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<5>.MM_i_24_1_48 XI0.XI1.XI3.XI3<5>.Y XI0.XI1.XI3.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<5>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<4>.MM_i_0 VSS! XI0.XI1.XI3.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<4>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<4>.MM_i_0_15 VSS! REG_DATA_12<4> XI0.XI1.XI3.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<4>.MM_i_0_15_63 XI0.XI1.XI3.XI3<4>.DUMMY1 REG_DATA_12<4>
+ XI0.XI1.XI3.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<4>.NEN
+ XI0.XI1.XI3.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<4>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<4>.MM_i_24 VDD! XI0.XI1.XI3.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<4>.MM_i_24_1 XI0.XI1.XI3.XI3<4>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<4>.MM_i_24_0 VDD! REG_DATA_12<4> XI0.XI1.XI3.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_12<4> XI0.XI1.XI3.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<4>.MM_i_24_1_48 XI0.XI1.XI3.XI3<4>.Y XI0.XI1.XI3.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<4>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<11>.MM_i_0 VSS! XI0.XI1.XI3.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<11>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<11>.MM_i_0_15 VSS! REG_DATA_12<11> XI0.XI1.XI3.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<11>.MM_i_0_15_63 XI0.XI1.XI3.XI3<11>.DUMMY1 REG_DATA_12<11>
+ XI0.XI1.XI3.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<11>.NEN
+ XI0.XI1.XI3.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<11>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<11>.MM_i_24 VDD! XI0.XI1.XI3.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<11>.MM_i_24_1 XI0.XI1.XI3.XI3<11>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<11>.MM_i_24_0 VDD! REG_DATA_12<11> XI0.XI1.XI3.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_12<11> XI0.XI1.XI3.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<11>.MM_i_24_1_48 XI0.XI1.XI3.XI3<11>.Y XI0.XI1.XI3.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<11>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<10>.MM_i_0 VSS! XI0.XI1.XI3.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<10>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<10>.MM_i_0_15 VSS! REG_DATA_12<10> XI0.XI1.XI3.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<10>.MM_i_0_15_63 XI0.XI1.XI3.XI3<10>.DUMMY1 REG_DATA_12<10>
+ XI0.XI1.XI3.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<10>.NEN
+ XI0.XI1.XI3.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<10>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<10>.MM_i_24 VDD! XI0.XI1.XI3.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<10>.MM_i_24_1 XI0.XI1.XI3.XI3<10>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<10>.MM_i_24_0 VDD! REG_DATA_12<10> XI0.XI1.XI3.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_12<10> XI0.XI1.XI3.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<10>.MM_i_24_1_48 XI0.XI1.XI3.XI3<10>.Y XI0.XI1.XI3.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<10>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<9>.MM_i_0 VSS! XI0.XI1.XI3.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<9>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<9>.MM_i_0_15 VSS! REG_DATA_12<9> XI0.XI1.XI3.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<9>.MM_i_0_15_63 XI0.XI1.XI3.XI3<9>.DUMMY1 REG_DATA_12<9>
+ XI0.XI1.XI3.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<9>.NEN
+ XI0.XI1.XI3.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<9>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<9>.MM_i_24 VDD! XI0.XI1.XI3.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<9>.MM_i_24_1 XI0.XI1.XI3.XI3<9>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<9>.MM_i_24_0 VDD! REG_DATA_12<9> XI0.XI1.XI3.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_12<9> XI0.XI1.XI3.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<9>.MM_i_24_1_48 XI0.XI1.XI3.XI3<9>.Y XI0.XI1.XI3.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<9>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<8>.MM_i_0 VSS! XI0.XI1.XI3.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<8>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<8>.MM_i_0_15 VSS! REG_DATA_12<8> XI0.XI1.XI3.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<8>.MM_i_0_15_63 XI0.XI1.XI3.XI3<8>.DUMMY1 REG_DATA_12<8>
+ XI0.XI1.XI3.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<8>.NEN
+ XI0.XI1.XI3.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<8>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<8>.MM_i_24 VDD! XI0.XI1.XI3.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<8>.MM_i_24_1 XI0.XI1.XI3.XI3<8>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<8>.MM_i_24_0 VDD! REG_DATA_12<8> XI0.XI1.XI3.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_12<8> XI0.XI1.XI3.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI3.XI3<8>.MM_i_24_1_48 XI0.XI1.XI3.XI3<8>.Y XI0.XI1.XI3.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<8>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<15>.MM_i_0 VSS! XI0.XI1.XI3.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<15>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<15>.MM_i_0_15 VSS! REG_DATA_12<15> XI0.XI1.XI3.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<15>.MM_i_0_15_63 XI0.XI1.XI3.XI3<15>.DUMMY1 REG_DATA_12<15>
+ XI0.XI1.XI3.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<15>.NEN
+ XI0.XI1.XI3.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<15>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<15>.MM_i_24 VDD! XI0.XI1.XI3.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<15>.MM_i_24_1 XI0.XI1.XI3.XI3<15>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<15>.MM_i_24_0 VDD! REG_DATA_12<15> XI0.XI1.XI3.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_12<15> XI0.XI1.XI3.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<15>.MM_i_24_1_48 XI0.XI1.XI3.XI3<15>.Y XI0.XI1.XI3.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<15>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<14>.MM_i_0 VSS! XI0.XI1.XI3.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<14>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<14>.MM_i_0_15 VSS! REG_DATA_12<14> XI0.XI1.XI3.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<14>.MM_i_0_15_63 XI0.XI1.XI3.XI3<14>.DUMMY1 REG_DATA_12<14>
+ XI0.XI1.XI3.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<14>.NEN
+ XI0.XI1.XI3.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<14>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<14>.MM_i_24 VDD! XI0.XI1.XI3.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<14>.MM_i_24_1 XI0.XI1.XI3.XI3<14>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<14>.MM_i_24_0 VDD! REG_DATA_12<14> XI0.XI1.XI3.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_12<14> XI0.XI1.XI3.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<14>.MM_i_24_1_48 XI0.XI1.XI3.XI3<14>.Y XI0.XI1.XI3.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<14>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<13>.MM_i_0 VSS! XI0.XI1.XI3.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<13>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<13>.MM_i_0_15 VSS! REG_DATA_12<13> XI0.XI1.XI3.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<13>.MM_i_0_15_63 XI0.XI1.XI3.XI3<13>.DUMMY1 REG_DATA_12<13>
+ XI0.XI1.XI3.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<13>.NEN
+ XI0.XI1.XI3.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<13>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<13>.MM_i_24 VDD! XI0.XI1.XI3.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<13>.MM_i_24_1 XI0.XI1.XI3.XI3<13>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<13>.MM_i_24_0 VDD! REG_DATA_12<13> XI0.XI1.XI3.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_12<13> XI0.XI1.XI3.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<13>.MM_i_24_1_48 XI0.XI1.XI3.XI3<13>.Y XI0.XI1.XI3.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<13>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI3.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI3.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI3.XI3<12>.MM_i_0 VSS! XI0.XI1.XI3.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI3.XI3<12>.MM_i_0_14 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<12>.MM_i_0_15 VSS! REG_DATA_12<12> XI0.XI1.XI3.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<12>.MM_i_0_15_63 XI0.XI1.XI3.XI3<12>.DUMMY1 REG_DATA_12<12>
+ XI0.XI1.XI3.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI3.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI3.XI3<12>.NEN
+ XI0.XI1.XI3.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI3.XI3<12>.MM_i_17 VSS! XI0.NET1<0> XI0.XI1.XI3.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI3.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI3.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<12>.MM_i_24 VDD! XI0.XI1.XI3.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI3.XI3<12>.MM_i_24_1 XI0.XI1.XI3.XI3<12>.DUMMY0 XI0.NET1<0>
+ XI0.XI1.XI3.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI3.XI3<12>.MM_i_24_0 VDD! REG_DATA_12<12> XI0.XI1.XI3.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_12<12> XI0.XI1.XI3.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI3.XI3<12>.MM_i_24_1_48 XI0.XI1.XI3.XI3<12>.Y XI0.XI1.XI3.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI3.XI3<12>.MM_i_42 VDD! XI0.NET1<0> XI0.XI1.XI3.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<3>.MM_i_0 VSS! XI0.XI1.XI4.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<3>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<3>.MM_i_0_15 VSS! REG_DATA_11<3> XI0.XI1.XI4.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<3>.MM_i_0_15_63 XI0.XI1.XI4.XI3<3>.DUMMY1 REG_DATA_11<3>
+ XI0.XI1.XI4.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<3>.NEN
+ XI0.XI1.XI4.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<3>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<3>.MM_i_24 VDD! XI0.XI1.XI4.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<3>.MM_i_24_1 XI0.XI1.XI4.XI3<3>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<3>.MM_i_24_0 VDD! REG_DATA_11<3> XI0.XI1.XI4.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_11<3> XI0.XI1.XI4.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<3>.MM_i_24_1_48 XI0.XI1.XI4.XI3<3>.Y XI0.XI1.XI4.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<3>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<2>.MM_i_0 VSS! XI0.XI1.XI4.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<2>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<2>.MM_i_0_15 VSS! REG_DATA_11<2> XI0.XI1.XI4.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<2>.MM_i_0_15_63 XI0.XI1.XI4.XI3<2>.DUMMY1 REG_DATA_11<2>
+ XI0.XI1.XI4.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<2>.NEN
+ XI0.XI1.XI4.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<2>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<2>.MM_i_24 VDD! XI0.XI1.XI4.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<2>.MM_i_24_1 XI0.XI1.XI4.XI3<2>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<2>.MM_i_24_0 VDD! REG_DATA_11<2> XI0.XI1.XI4.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_11<2> XI0.XI1.XI4.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<2>.MM_i_24_1_48 XI0.XI1.XI4.XI3<2>.Y XI0.XI1.XI4.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<2>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<1>.MM_i_0 VSS! XI0.XI1.XI4.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<1>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<1>.MM_i_0_15 VSS! REG_DATA_11<1> XI0.XI1.XI4.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<1>.MM_i_0_15_63 XI0.XI1.XI4.XI3<1>.DUMMY1 REG_DATA_11<1>
+ XI0.XI1.XI4.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<1>.NEN
+ XI0.XI1.XI4.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<1>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<1>.MM_i_24 VDD! XI0.XI1.XI4.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<1>.MM_i_24_1 XI0.XI1.XI4.XI3<1>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<1>.MM_i_24_0 VDD! REG_DATA_11<1> XI0.XI1.XI4.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_11<1> XI0.XI1.XI4.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<1>.MM_i_24_1_48 XI0.XI1.XI4.XI3<1>.Y XI0.XI1.XI4.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<1>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<0>.MM_i_0 VSS! XI0.XI1.XI4.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<0>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<0>.MM_i_0_15 VSS! REG_DATA_11<0> XI0.XI1.XI4.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<0>.MM_i_0_15_63 XI0.XI1.XI4.XI3<0>.DUMMY1 REG_DATA_11<0>
+ XI0.XI1.XI4.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<0>.NEN
+ XI0.XI1.XI4.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<0>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<0>.MM_i_24 VDD! XI0.XI1.XI4.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<0>.MM_i_24_1 XI0.XI1.XI4.XI3<0>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<0>.MM_i_24_0 VDD! REG_DATA_11<0> XI0.XI1.XI4.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_11<0> XI0.XI1.XI4.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<0>.MM_i_24_1_48 XI0.XI1.XI4.XI3<0>.Y XI0.XI1.XI4.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<0>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<7>.MM_i_0 VSS! XI0.XI1.XI4.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<7>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<7>.MM_i_0_15 VSS! REG_DATA_11<7> XI0.XI1.XI4.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<7>.MM_i_0_15_63 XI0.XI1.XI4.XI3<7>.DUMMY1 REG_DATA_11<7>
+ XI0.XI1.XI4.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<7>.NEN
+ XI0.XI1.XI4.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<7>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<7>.MM_i_24 VDD! XI0.XI1.XI4.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<7>.MM_i_24_1 XI0.XI1.XI4.XI3<7>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<7>.MM_i_24_0 VDD! REG_DATA_11<7> XI0.XI1.XI4.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_11<7> XI0.XI1.XI4.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<7>.MM_i_24_1_48 XI0.XI1.XI4.XI3<7>.Y XI0.XI1.XI4.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<7>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<6>.MM_i_0 VSS! XI0.XI1.XI4.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<6>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<6>.MM_i_0_15 VSS! REG_DATA_11<6> XI0.XI1.XI4.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<6>.MM_i_0_15_63 XI0.XI1.XI4.XI3<6>.DUMMY1 REG_DATA_11<6>
+ XI0.XI1.XI4.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<6>.NEN
+ XI0.XI1.XI4.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<6>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<6>.MM_i_24 VDD! XI0.XI1.XI4.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<6>.MM_i_24_1 XI0.XI1.XI4.XI3<6>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<6>.MM_i_24_0 VDD! REG_DATA_11<6> XI0.XI1.XI4.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_11<6> XI0.XI1.XI4.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<6>.MM_i_24_1_48 XI0.XI1.XI4.XI3<6>.Y XI0.XI1.XI4.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<6>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<5>.MM_i_0 VSS! XI0.XI1.XI4.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<5>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<5>.MM_i_0_15 VSS! REG_DATA_11<5> XI0.XI1.XI4.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<5>.MM_i_0_15_63 XI0.XI1.XI4.XI3<5>.DUMMY1 REG_DATA_11<5>
+ XI0.XI1.XI4.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<5>.NEN
+ XI0.XI1.XI4.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<5>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<5>.MM_i_24 VDD! XI0.XI1.XI4.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<5>.MM_i_24_1 XI0.XI1.XI4.XI3<5>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<5>.MM_i_24_0 VDD! REG_DATA_11<5> XI0.XI1.XI4.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_11<5> XI0.XI1.XI4.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<5>.MM_i_24_1_48 XI0.XI1.XI4.XI3<5>.Y XI0.XI1.XI4.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<5>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<4>.MM_i_0 VSS! XI0.XI1.XI4.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<4>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<4>.MM_i_0_15 VSS! REG_DATA_11<4> XI0.XI1.XI4.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<4>.MM_i_0_15_63 XI0.XI1.XI4.XI3<4>.DUMMY1 REG_DATA_11<4>
+ XI0.XI1.XI4.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<4>.NEN
+ XI0.XI1.XI4.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<4>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<4>.MM_i_24 VDD! XI0.XI1.XI4.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<4>.MM_i_24_1 XI0.XI1.XI4.XI3<4>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<4>.MM_i_24_0 VDD! REG_DATA_11<4> XI0.XI1.XI4.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_11<4> XI0.XI1.XI4.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<4>.MM_i_24_1_48 XI0.XI1.XI4.XI3<4>.Y XI0.XI1.XI4.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<4>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<11>.MM_i_0 VSS! XI0.XI1.XI4.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<11>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<11>.MM_i_0_15 VSS! REG_DATA_11<11> XI0.XI1.XI4.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<11>.MM_i_0_15_63 XI0.XI1.XI4.XI3<11>.DUMMY1 REG_DATA_11<11>
+ XI0.XI1.XI4.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<11>.NEN
+ XI0.XI1.XI4.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<11>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<11>.MM_i_24 VDD! XI0.XI1.XI4.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<11>.MM_i_24_1 XI0.XI1.XI4.XI3<11>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<11>.MM_i_24_0 VDD! REG_DATA_11<11> XI0.XI1.XI4.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_11<11> XI0.XI1.XI4.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<11>.MM_i_24_1_48 XI0.XI1.XI4.XI3<11>.Y XI0.XI1.XI4.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<11>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<10>.MM_i_0 VSS! XI0.XI1.XI4.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<10>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<10>.MM_i_0_15 VSS! REG_DATA_11<10> XI0.XI1.XI4.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<10>.MM_i_0_15_63 XI0.XI1.XI4.XI3<10>.DUMMY1 REG_DATA_11<10>
+ XI0.XI1.XI4.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<10>.NEN
+ XI0.XI1.XI4.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<10>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<10>.MM_i_24 VDD! XI0.XI1.XI4.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<10>.MM_i_24_1 XI0.XI1.XI4.XI3<10>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<10>.MM_i_24_0 VDD! REG_DATA_11<10> XI0.XI1.XI4.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_11<10> XI0.XI1.XI4.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<10>.MM_i_24_1_48 XI0.XI1.XI4.XI3<10>.Y XI0.XI1.XI4.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<10>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<9>.MM_i_0 VSS! XI0.XI1.XI4.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<9>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<9>.MM_i_0_15 VSS! REG_DATA_11<9> XI0.XI1.XI4.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<9>.MM_i_0_15_63 XI0.XI1.XI4.XI3<9>.DUMMY1 REG_DATA_11<9>
+ XI0.XI1.XI4.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<9>.NEN
+ XI0.XI1.XI4.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<9>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<9>.MM_i_24 VDD! XI0.XI1.XI4.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<9>.MM_i_24_1 XI0.XI1.XI4.XI3<9>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<9>.MM_i_24_0 VDD! REG_DATA_11<9> XI0.XI1.XI4.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_11<9> XI0.XI1.XI4.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<9>.MM_i_24_1_48 XI0.XI1.XI4.XI3<9>.Y XI0.XI1.XI4.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<9>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<8>.MM_i_0 VSS! XI0.XI1.XI4.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<8>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<8>.MM_i_0_15 VSS! REG_DATA_11<8> XI0.XI1.XI4.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<8>.MM_i_0_15_63 XI0.XI1.XI4.XI3<8>.DUMMY1 REG_DATA_11<8>
+ XI0.XI1.XI4.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<8>.NEN
+ XI0.XI1.XI4.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<8>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<8>.MM_i_24 VDD! XI0.XI1.XI4.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<8>.MM_i_24_1 XI0.XI1.XI4.XI3<8>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<8>.MM_i_24_0 VDD! REG_DATA_11<8> XI0.XI1.XI4.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_11<8> XI0.XI1.XI4.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI4.XI3<8>.MM_i_24_1_48 XI0.XI1.XI4.XI3<8>.Y XI0.XI1.XI4.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<8>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<15>.MM_i_0 VSS! XI0.XI1.XI4.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<15>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<15>.MM_i_0_15 VSS! REG_DATA_11<15> XI0.XI1.XI4.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<15>.MM_i_0_15_63 XI0.XI1.XI4.XI3<15>.DUMMY1 REG_DATA_11<15>
+ XI0.XI1.XI4.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<15>.NEN
+ XI0.XI1.XI4.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<15>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<15>.MM_i_24 VDD! XI0.XI1.XI4.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<15>.MM_i_24_1 XI0.XI1.XI4.XI3<15>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<15>.MM_i_24_0 VDD! REG_DATA_11<15> XI0.XI1.XI4.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_11<15> XI0.XI1.XI4.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<15>.MM_i_24_1_48 XI0.XI1.XI4.XI3<15>.Y XI0.XI1.XI4.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<15>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<14>.MM_i_0 VSS! XI0.XI1.XI4.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<14>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<14>.MM_i_0_15 VSS! REG_DATA_11<14> XI0.XI1.XI4.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<14>.MM_i_0_15_63 XI0.XI1.XI4.XI3<14>.DUMMY1 REG_DATA_11<14>
+ XI0.XI1.XI4.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<14>.NEN
+ XI0.XI1.XI4.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<14>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<14>.MM_i_24 VDD! XI0.XI1.XI4.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<14>.MM_i_24_1 XI0.XI1.XI4.XI3<14>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<14>.MM_i_24_0 VDD! REG_DATA_11<14> XI0.XI1.XI4.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_11<14> XI0.XI1.XI4.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<14>.MM_i_24_1_48 XI0.XI1.XI4.XI3<14>.Y XI0.XI1.XI4.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<14>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<13>.MM_i_0 VSS! XI0.XI1.XI4.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<13>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<13>.MM_i_0_15 VSS! REG_DATA_11<13> XI0.XI1.XI4.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<13>.MM_i_0_15_63 XI0.XI1.XI4.XI3<13>.DUMMY1 REG_DATA_11<13>
+ XI0.XI1.XI4.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<13>.NEN
+ XI0.XI1.XI4.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<13>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<13>.MM_i_24 VDD! XI0.XI1.XI4.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<13>.MM_i_24_1 XI0.XI1.XI4.XI3<13>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<13>.MM_i_24_0 VDD! REG_DATA_11<13> XI0.XI1.XI4.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_11<13> XI0.XI1.XI4.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<13>.MM_i_24_1_48 XI0.XI1.XI4.XI3<13>.Y XI0.XI1.XI4.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<13>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI4.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI4.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI4.XI3<12>.MM_i_0 VSS! XI0.XI1.XI4.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI4.XI3<12>.MM_i_0_14 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<12>.MM_i_0_15 VSS! REG_DATA_11<12> XI0.XI1.XI4.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<12>.MM_i_0_15_63 XI0.XI1.XI4.XI3<12>.DUMMY1 REG_DATA_11<12>
+ XI0.XI1.XI4.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI4.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI4.XI3<12>.NEN
+ XI0.XI1.XI4.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI4.XI3<12>.MM_i_17 VSS! XI0.NET1<1> XI0.XI1.XI4.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI4.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI4.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<12>.MM_i_24 VDD! XI0.XI1.XI4.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI4.XI3<12>.MM_i_24_1 XI0.XI1.XI4.XI3<12>.DUMMY0 XI0.NET1<1>
+ XI0.XI1.XI4.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI4.XI3<12>.MM_i_24_0 VDD! REG_DATA_11<12> XI0.XI1.XI4.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_11<12> XI0.XI1.XI4.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI4.XI3<12>.MM_i_24_1_48 XI0.XI1.XI4.XI3<12>.Y XI0.XI1.XI4.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI4.XI3<12>.MM_i_42 VDD! XI0.NET1<1> XI0.XI1.XI4.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<3>.MM_i_0 VSS! XI0.XI1.XI6.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<3>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<3>.MM_i_0_15 VSS! REG_DATA_10<3> XI0.XI1.XI6.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<3>.MM_i_0_15_63 XI0.XI1.XI6.XI3<3>.DUMMY1 REG_DATA_10<3>
+ XI0.XI1.XI6.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<3>.NEN
+ XI0.XI1.XI6.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<3>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<3>.MM_i_24 VDD! XI0.XI1.XI6.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<3>.MM_i_24_1 XI0.XI1.XI6.XI3<3>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<3>.MM_i_24_0 VDD! REG_DATA_10<3> XI0.XI1.XI6.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_10<3> XI0.XI1.XI6.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<3>.MM_i_24_1_48 XI0.XI1.XI6.XI3<3>.Y XI0.XI1.XI6.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<3>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<2>.MM_i_0 VSS! XI0.XI1.XI6.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<2>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<2>.MM_i_0_15 VSS! REG_DATA_10<2> XI0.XI1.XI6.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<2>.MM_i_0_15_63 XI0.XI1.XI6.XI3<2>.DUMMY1 REG_DATA_10<2>
+ XI0.XI1.XI6.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<2>.NEN
+ XI0.XI1.XI6.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<2>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<2>.MM_i_24 VDD! XI0.XI1.XI6.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<2>.MM_i_24_1 XI0.XI1.XI6.XI3<2>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<2>.MM_i_24_0 VDD! REG_DATA_10<2> XI0.XI1.XI6.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_10<2> XI0.XI1.XI6.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<2>.MM_i_24_1_48 XI0.XI1.XI6.XI3<2>.Y XI0.XI1.XI6.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<2>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<1>.MM_i_0 VSS! XI0.XI1.XI6.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<1>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<1>.MM_i_0_15 VSS! REG_DATA_10<1> XI0.XI1.XI6.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<1>.MM_i_0_15_63 XI0.XI1.XI6.XI3<1>.DUMMY1 REG_DATA_10<1>
+ XI0.XI1.XI6.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<1>.NEN
+ XI0.XI1.XI6.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<1>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<1>.MM_i_24 VDD! XI0.XI1.XI6.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<1>.MM_i_24_1 XI0.XI1.XI6.XI3<1>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<1>.MM_i_24_0 VDD! REG_DATA_10<1> XI0.XI1.XI6.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_10<1> XI0.XI1.XI6.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<1>.MM_i_24_1_48 XI0.XI1.XI6.XI3<1>.Y XI0.XI1.XI6.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<1>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<0>.MM_i_0 VSS! XI0.XI1.XI6.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<0>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<0>.MM_i_0_15 VSS! REG_DATA_10<0> XI0.XI1.XI6.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<0>.MM_i_0_15_63 XI0.XI1.XI6.XI3<0>.DUMMY1 REG_DATA_10<0>
+ XI0.XI1.XI6.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<0>.NEN
+ XI0.XI1.XI6.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<0>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<0>.MM_i_24 VDD! XI0.XI1.XI6.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<0>.MM_i_24_1 XI0.XI1.XI6.XI3<0>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<0>.MM_i_24_0 VDD! REG_DATA_10<0> XI0.XI1.XI6.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_10<0> XI0.XI1.XI6.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<0>.MM_i_24_1_48 XI0.XI1.XI6.XI3<0>.Y XI0.XI1.XI6.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<0>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<7>.MM_i_0 VSS! XI0.XI1.XI6.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<7>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<7>.MM_i_0_15 VSS! REG_DATA_10<7> XI0.XI1.XI6.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<7>.MM_i_0_15_63 XI0.XI1.XI6.XI3<7>.DUMMY1 REG_DATA_10<7>
+ XI0.XI1.XI6.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<7>.NEN
+ XI0.XI1.XI6.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<7>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<7>.MM_i_24 VDD! XI0.XI1.XI6.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<7>.MM_i_24_1 XI0.XI1.XI6.XI3<7>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<7>.MM_i_24_0 VDD! REG_DATA_10<7> XI0.XI1.XI6.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_10<7> XI0.XI1.XI6.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<7>.MM_i_24_1_48 XI0.XI1.XI6.XI3<7>.Y XI0.XI1.XI6.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<7>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<6>.MM_i_0 VSS! XI0.XI1.XI6.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<6>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<6>.MM_i_0_15 VSS! REG_DATA_10<6> XI0.XI1.XI6.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<6>.MM_i_0_15_63 XI0.XI1.XI6.XI3<6>.DUMMY1 REG_DATA_10<6>
+ XI0.XI1.XI6.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<6>.NEN
+ XI0.XI1.XI6.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<6>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<6>.MM_i_24 VDD! XI0.XI1.XI6.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<6>.MM_i_24_1 XI0.XI1.XI6.XI3<6>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<6>.MM_i_24_0 VDD! REG_DATA_10<6> XI0.XI1.XI6.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_10<6> XI0.XI1.XI6.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<6>.MM_i_24_1_48 XI0.XI1.XI6.XI3<6>.Y XI0.XI1.XI6.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<6>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<5>.MM_i_0 VSS! XI0.XI1.XI6.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<5>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<5>.MM_i_0_15 VSS! REG_DATA_10<5> XI0.XI1.XI6.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<5>.MM_i_0_15_63 XI0.XI1.XI6.XI3<5>.DUMMY1 REG_DATA_10<5>
+ XI0.XI1.XI6.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<5>.NEN
+ XI0.XI1.XI6.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<5>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<5>.MM_i_24 VDD! XI0.XI1.XI6.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<5>.MM_i_24_1 XI0.XI1.XI6.XI3<5>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<5>.MM_i_24_0 VDD! REG_DATA_10<5> XI0.XI1.XI6.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_10<5> XI0.XI1.XI6.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<5>.MM_i_24_1_48 XI0.XI1.XI6.XI3<5>.Y XI0.XI1.XI6.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<5>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<4>.MM_i_0 VSS! XI0.XI1.XI6.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<4>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<4>.MM_i_0_15 VSS! REG_DATA_10<4> XI0.XI1.XI6.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<4>.MM_i_0_15_63 XI0.XI1.XI6.XI3<4>.DUMMY1 REG_DATA_10<4>
+ XI0.XI1.XI6.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<4>.NEN
+ XI0.XI1.XI6.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<4>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<4>.MM_i_24 VDD! XI0.XI1.XI6.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<4>.MM_i_24_1 XI0.XI1.XI6.XI3<4>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<4>.MM_i_24_0 VDD! REG_DATA_10<4> XI0.XI1.XI6.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_10<4> XI0.XI1.XI6.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<4>.MM_i_24_1_48 XI0.XI1.XI6.XI3<4>.Y XI0.XI1.XI6.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<4>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<11>.MM_i_0 VSS! XI0.XI1.XI6.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<11>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<11>.MM_i_0_15 VSS! REG_DATA_10<11> XI0.XI1.XI6.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<11>.MM_i_0_15_63 XI0.XI1.XI6.XI3<11>.DUMMY1 REG_DATA_10<11>
+ XI0.XI1.XI6.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<11>.NEN
+ XI0.XI1.XI6.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<11>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<11>.MM_i_24 VDD! XI0.XI1.XI6.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<11>.MM_i_24_1 XI0.XI1.XI6.XI3<11>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<11>.MM_i_24_0 VDD! REG_DATA_10<11> XI0.XI1.XI6.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_10<11> XI0.XI1.XI6.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<11>.MM_i_24_1_48 XI0.XI1.XI6.XI3<11>.Y XI0.XI1.XI6.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<11>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<10>.MM_i_0 VSS! XI0.XI1.XI6.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<10>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<10>.MM_i_0_15 VSS! REG_DATA_10<10> XI0.XI1.XI6.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<10>.MM_i_0_15_63 XI0.XI1.XI6.XI3<10>.DUMMY1 REG_DATA_10<10>
+ XI0.XI1.XI6.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<10>.NEN
+ XI0.XI1.XI6.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<10>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<10>.MM_i_24 VDD! XI0.XI1.XI6.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<10>.MM_i_24_1 XI0.XI1.XI6.XI3<10>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<10>.MM_i_24_0 VDD! REG_DATA_10<10> XI0.XI1.XI6.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_10<10> XI0.XI1.XI6.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<10>.MM_i_24_1_48 XI0.XI1.XI6.XI3<10>.Y XI0.XI1.XI6.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<10>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<9>.MM_i_0 VSS! XI0.XI1.XI6.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<9>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<9>.MM_i_0_15 VSS! REG_DATA_10<9> XI0.XI1.XI6.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<9>.MM_i_0_15_63 XI0.XI1.XI6.XI3<9>.DUMMY1 REG_DATA_10<9>
+ XI0.XI1.XI6.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<9>.NEN
+ XI0.XI1.XI6.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<9>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<9>.MM_i_24 VDD! XI0.XI1.XI6.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<9>.MM_i_24_1 XI0.XI1.XI6.XI3<9>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<9>.MM_i_24_0 VDD! REG_DATA_10<9> XI0.XI1.XI6.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_10<9> XI0.XI1.XI6.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<9>.MM_i_24_1_48 XI0.XI1.XI6.XI3<9>.Y XI0.XI1.XI6.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<9>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<8>.MM_i_0 VSS! XI0.XI1.XI6.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<8>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<8>.MM_i_0_15 VSS! REG_DATA_10<8> XI0.XI1.XI6.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<8>.MM_i_0_15_63 XI0.XI1.XI6.XI3<8>.DUMMY1 REG_DATA_10<8>
+ XI0.XI1.XI6.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<8>.NEN
+ XI0.XI1.XI6.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<8>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<8>.MM_i_24 VDD! XI0.XI1.XI6.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<8>.MM_i_24_1 XI0.XI1.XI6.XI3<8>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<8>.MM_i_24_0 VDD! REG_DATA_10<8> XI0.XI1.XI6.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_10<8> XI0.XI1.XI6.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI6.XI3<8>.MM_i_24_1_48 XI0.XI1.XI6.XI3<8>.Y XI0.XI1.XI6.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<8>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<15>.MM_i_0 VSS! XI0.XI1.XI6.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<15>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<15>.MM_i_0_15 VSS! REG_DATA_10<15> XI0.XI1.XI6.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<15>.MM_i_0_15_63 XI0.XI1.XI6.XI3<15>.DUMMY1 REG_DATA_10<15>
+ XI0.XI1.XI6.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<15>.NEN
+ XI0.XI1.XI6.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<15>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<15>.MM_i_24 VDD! XI0.XI1.XI6.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<15>.MM_i_24_1 XI0.XI1.XI6.XI3<15>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<15>.MM_i_24_0 VDD! REG_DATA_10<15> XI0.XI1.XI6.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_10<15> XI0.XI1.XI6.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<15>.MM_i_24_1_48 XI0.XI1.XI6.XI3<15>.Y XI0.XI1.XI6.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<15>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<14>.MM_i_0 VSS! XI0.XI1.XI6.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<14>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<14>.MM_i_0_15 VSS! REG_DATA_10<14> XI0.XI1.XI6.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<14>.MM_i_0_15_63 XI0.XI1.XI6.XI3<14>.DUMMY1 REG_DATA_10<14>
+ XI0.XI1.XI6.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<14>.NEN
+ XI0.XI1.XI6.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<14>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<14>.MM_i_24 VDD! XI0.XI1.XI6.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<14>.MM_i_24_1 XI0.XI1.XI6.XI3<14>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<14>.MM_i_24_0 VDD! REG_DATA_10<14> XI0.XI1.XI6.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_10<14> XI0.XI1.XI6.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<14>.MM_i_24_1_48 XI0.XI1.XI6.XI3<14>.Y XI0.XI1.XI6.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<14>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<13>.MM_i_0 VSS! XI0.XI1.XI6.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<13>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<13>.MM_i_0_15 VSS! REG_DATA_10<13> XI0.XI1.XI6.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<13>.MM_i_0_15_63 XI0.XI1.XI6.XI3<13>.DUMMY1 REG_DATA_10<13>
+ XI0.XI1.XI6.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<13>.NEN
+ XI0.XI1.XI6.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<13>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<13>.MM_i_24 VDD! XI0.XI1.XI6.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<13>.MM_i_24_1 XI0.XI1.XI6.XI3<13>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<13>.MM_i_24_0 VDD! REG_DATA_10<13> XI0.XI1.XI6.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_10<13> XI0.XI1.XI6.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<13>.MM_i_24_1_48 XI0.XI1.XI6.XI3<13>.Y XI0.XI1.XI6.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<13>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI6.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI6.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI6.XI3<12>.MM_i_0 VSS! XI0.XI1.XI6.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI6.XI3<12>.MM_i_0_14 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<12>.MM_i_0_15 VSS! REG_DATA_10<12> XI0.XI1.XI6.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<12>.MM_i_0_15_63 XI0.XI1.XI6.XI3<12>.DUMMY1 REG_DATA_10<12>
+ XI0.XI1.XI6.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI6.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI6.XI3<12>.NEN
+ XI0.XI1.XI6.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI6.XI3<12>.MM_i_17 VSS! XI0.NET1<2> XI0.XI1.XI6.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI6.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI6.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<12>.MM_i_24 VDD! XI0.XI1.XI6.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI6.XI3<12>.MM_i_24_1 XI0.XI1.XI6.XI3<12>.DUMMY0 XI0.NET1<2>
+ XI0.XI1.XI6.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI6.XI3<12>.MM_i_24_0 VDD! REG_DATA_10<12> XI0.XI1.XI6.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_10<12> XI0.XI1.XI6.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI6.XI3<12>.MM_i_24_1_48 XI0.XI1.XI6.XI3<12>.Y XI0.XI1.XI6.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI6.XI3<12>.MM_i_42 VDD! XI0.NET1<2> XI0.XI1.XI6.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<3>.MM_i_0 VSS! XI0.XI1.XI5.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<3>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<3>.MM_i_0_15 VSS! REG_DATA_9<3> XI0.XI1.XI5.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<3>.MM_i_0_15_63 XI0.XI1.XI5.XI3<3>.DUMMY1 REG_DATA_9<3>
+ XI0.XI1.XI5.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<3>.NEN
+ XI0.XI1.XI5.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<3>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<3>.MM_i_24 VDD! XI0.XI1.XI5.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<3>.MM_i_24_1 XI0.XI1.XI5.XI3<3>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<3>.MM_i_24_0 VDD! REG_DATA_9<3> XI0.XI1.XI5.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_9<3> XI0.XI1.XI5.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<3>.MM_i_24_1_48 XI0.XI1.XI5.XI3<3>.Y XI0.XI1.XI5.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<3>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<2>.MM_i_0 VSS! XI0.XI1.XI5.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<2>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<2>.MM_i_0_15 VSS! REG_DATA_9<2> XI0.XI1.XI5.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<2>.MM_i_0_15_63 XI0.XI1.XI5.XI3<2>.DUMMY1 REG_DATA_9<2>
+ XI0.XI1.XI5.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<2>.NEN
+ XI0.XI1.XI5.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<2>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<2>.MM_i_24 VDD! XI0.XI1.XI5.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<2>.MM_i_24_1 XI0.XI1.XI5.XI3<2>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<2>.MM_i_24_0 VDD! REG_DATA_9<2> XI0.XI1.XI5.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_9<2> XI0.XI1.XI5.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<2>.MM_i_24_1_48 XI0.XI1.XI5.XI3<2>.Y XI0.XI1.XI5.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<2>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<1>.MM_i_0 VSS! XI0.XI1.XI5.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<1>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<1>.MM_i_0_15 VSS! REG_DATA_9<1> XI0.XI1.XI5.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<1>.MM_i_0_15_63 XI0.XI1.XI5.XI3<1>.DUMMY1 REG_DATA_9<1>
+ XI0.XI1.XI5.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<1>.NEN
+ XI0.XI1.XI5.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<1>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<1>.MM_i_24 VDD! XI0.XI1.XI5.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<1>.MM_i_24_1 XI0.XI1.XI5.XI3<1>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<1>.MM_i_24_0 VDD! REG_DATA_9<1> XI0.XI1.XI5.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_9<1> XI0.XI1.XI5.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<1>.MM_i_24_1_48 XI0.XI1.XI5.XI3<1>.Y XI0.XI1.XI5.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<1>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<0>.MM_i_0 VSS! XI0.XI1.XI5.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<0>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<0>.MM_i_0_15 VSS! REG_DATA_9<0> XI0.XI1.XI5.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<0>.MM_i_0_15_63 XI0.XI1.XI5.XI3<0>.DUMMY1 REG_DATA_9<0>
+ XI0.XI1.XI5.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<0>.NEN
+ XI0.XI1.XI5.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<0>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<0>.MM_i_24 VDD! XI0.XI1.XI5.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<0>.MM_i_24_1 XI0.XI1.XI5.XI3<0>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<0>.MM_i_24_0 VDD! REG_DATA_9<0> XI0.XI1.XI5.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_9<0> XI0.XI1.XI5.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<0>.MM_i_24_1_48 XI0.XI1.XI5.XI3<0>.Y XI0.XI1.XI5.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<0>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<7>.MM_i_0 VSS! XI0.XI1.XI5.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<7>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<7>.MM_i_0_15 VSS! REG_DATA_9<7> XI0.XI1.XI5.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<7>.MM_i_0_15_63 XI0.XI1.XI5.XI3<7>.DUMMY1 REG_DATA_9<7>
+ XI0.XI1.XI5.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<7>.NEN
+ XI0.XI1.XI5.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<7>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<7>.MM_i_24 VDD! XI0.XI1.XI5.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<7>.MM_i_24_1 XI0.XI1.XI5.XI3<7>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<7>.MM_i_24_0 VDD! REG_DATA_9<7> XI0.XI1.XI5.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_9<7> XI0.XI1.XI5.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<7>.MM_i_24_1_48 XI0.XI1.XI5.XI3<7>.Y XI0.XI1.XI5.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<7>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<6>.MM_i_0 VSS! XI0.XI1.XI5.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<6>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<6>.MM_i_0_15 VSS! REG_DATA_9<6> XI0.XI1.XI5.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<6>.MM_i_0_15_63 XI0.XI1.XI5.XI3<6>.DUMMY1 REG_DATA_9<6>
+ XI0.XI1.XI5.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<6>.NEN
+ XI0.XI1.XI5.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<6>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<6>.MM_i_24 VDD! XI0.XI1.XI5.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<6>.MM_i_24_1 XI0.XI1.XI5.XI3<6>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<6>.MM_i_24_0 VDD! REG_DATA_9<6> XI0.XI1.XI5.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_9<6> XI0.XI1.XI5.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<6>.MM_i_24_1_48 XI0.XI1.XI5.XI3<6>.Y XI0.XI1.XI5.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<6>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<5>.MM_i_0 VSS! XI0.XI1.XI5.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<5>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<5>.MM_i_0_15 VSS! REG_DATA_9<5> XI0.XI1.XI5.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<5>.MM_i_0_15_63 XI0.XI1.XI5.XI3<5>.DUMMY1 REG_DATA_9<5>
+ XI0.XI1.XI5.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<5>.NEN
+ XI0.XI1.XI5.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<5>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<5>.MM_i_24 VDD! XI0.XI1.XI5.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<5>.MM_i_24_1 XI0.XI1.XI5.XI3<5>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<5>.MM_i_24_0 VDD! REG_DATA_9<5> XI0.XI1.XI5.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_9<5> XI0.XI1.XI5.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<5>.MM_i_24_1_48 XI0.XI1.XI5.XI3<5>.Y XI0.XI1.XI5.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<5>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<4>.MM_i_0 VSS! XI0.XI1.XI5.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<4>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<4>.MM_i_0_15 VSS! REG_DATA_9<4> XI0.XI1.XI5.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<4>.MM_i_0_15_63 XI0.XI1.XI5.XI3<4>.DUMMY1 REG_DATA_9<4>
+ XI0.XI1.XI5.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<4>.NEN
+ XI0.XI1.XI5.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<4>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<4>.MM_i_24 VDD! XI0.XI1.XI5.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<4>.MM_i_24_1 XI0.XI1.XI5.XI3<4>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<4>.MM_i_24_0 VDD! REG_DATA_9<4> XI0.XI1.XI5.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_9<4> XI0.XI1.XI5.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<4>.MM_i_24_1_48 XI0.XI1.XI5.XI3<4>.Y XI0.XI1.XI5.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<4>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<11>.MM_i_0 VSS! XI0.XI1.XI5.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<11>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<11>.MM_i_0_15 VSS! REG_DATA_9<11> XI0.XI1.XI5.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<11>.MM_i_0_15_63 XI0.XI1.XI5.XI3<11>.DUMMY1 REG_DATA_9<11>
+ XI0.XI1.XI5.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<11>.NEN
+ XI0.XI1.XI5.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<11>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<11>.MM_i_24 VDD! XI0.XI1.XI5.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<11>.MM_i_24_1 XI0.XI1.XI5.XI3<11>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<11>.MM_i_24_0 VDD! REG_DATA_9<11> XI0.XI1.XI5.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI5.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_9<11> XI0.XI1.XI5.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<11>.MM_i_24_1_48 XI0.XI1.XI5.XI3<11>.Y XI0.XI1.XI5.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<11>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<10>.MM_i_0 VSS! XI0.XI1.XI5.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<10>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<10>.MM_i_0_15 VSS! REG_DATA_9<10> XI0.XI1.XI5.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<10>.MM_i_0_15_63 XI0.XI1.XI5.XI3<10>.DUMMY1 REG_DATA_9<10>
+ XI0.XI1.XI5.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<10>.NEN
+ XI0.XI1.XI5.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<10>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<10>.MM_i_24 VDD! XI0.XI1.XI5.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<10>.MM_i_24_1 XI0.XI1.XI5.XI3<10>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<10>.MM_i_24_0 VDD! REG_DATA_9<10> XI0.XI1.XI5.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI5.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_9<10> XI0.XI1.XI5.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<10>.MM_i_24_1_48 XI0.XI1.XI5.XI3<10>.Y XI0.XI1.XI5.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<10>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<9>.MM_i_0 VSS! XI0.XI1.XI5.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<9>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<9>.MM_i_0_15 VSS! REG_DATA_9<9> XI0.XI1.XI5.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<9>.MM_i_0_15_63 XI0.XI1.XI5.XI3<9>.DUMMY1 REG_DATA_9<9>
+ XI0.XI1.XI5.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<9>.NEN
+ XI0.XI1.XI5.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<9>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<9>.MM_i_24 VDD! XI0.XI1.XI5.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<9>.MM_i_24_1 XI0.XI1.XI5.XI3<9>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<9>.MM_i_24_0 VDD! REG_DATA_9<9> XI0.XI1.XI5.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_9<9> XI0.XI1.XI5.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<9>.MM_i_24_1_48 XI0.XI1.XI5.XI3<9>.Y XI0.XI1.XI5.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<9>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<8>.MM_i_0 VSS! XI0.XI1.XI5.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<8>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<8>.MM_i_0_15 VSS! REG_DATA_9<8> XI0.XI1.XI5.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<8>.MM_i_0_15_63 XI0.XI1.XI5.XI3<8>.DUMMY1 REG_DATA_9<8>
+ XI0.XI1.XI5.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<8>.NEN
+ XI0.XI1.XI5.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<8>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<8>.MM_i_24 VDD! XI0.XI1.XI5.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<8>.MM_i_24_1 XI0.XI1.XI5.XI3<8>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<8>.MM_i_24_0 VDD! REG_DATA_9<8> XI0.XI1.XI5.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_9<8> XI0.XI1.XI5.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<8>.MM_i_24_1_48 XI0.XI1.XI5.XI3<8>.Y XI0.XI1.XI5.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<8>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<15>.MM_i_0 VSS! XI0.XI1.XI5.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<15>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<15>.MM_i_0_15 VSS! REG_DATA_9<15> XI0.XI1.XI5.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<15>.MM_i_0_15_63 XI0.XI1.XI5.XI3<15>.DUMMY1 REG_DATA_9<15>
+ XI0.XI1.XI5.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<15>.NEN
+ XI0.XI1.XI5.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<15>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<15>.MM_i_24 VDD! XI0.XI1.XI5.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<15>.MM_i_24_1 XI0.XI1.XI5.XI3<15>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<15>.MM_i_24_0 VDD! REG_DATA_9<15> XI0.XI1.XI5.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI5.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_9<15> XI0.XI1.XI5.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<15>.MM_i_24_1_48 XI0.XI1.XI5.XI3<15>.Y XI0.XI1.XI5.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<15>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<14>.MM_i_0 VSS! XI0.XI1.XI5.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<14>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<14>.MM_i_0_15 VSS! REG_DATA_9<14> XI0.XI1.XI5.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<14>.MM_i_0_15_63 XI0.XI1.XI5.XI3<14>.DUMMY1 REG_DATA_9<14>
+ XI0.XI1.XI5.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<14>.NEN
+ XI0.XI1.XI5.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<14>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<14>.MM_i_24 VDD! XI0.XI1.XI5.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<14>.MM_i_24_1 XI0.XI1.XI5.XI3<14>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<14>.MM_i_24_0 VDD! REG_DATA_9<14> XI0.XI1.XI5.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI5.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_9<14> XI0.XI1.XI5.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<14>.MM_i_24_1_48 XI0.XI1.XI5.XI3<14>.Y XI0.XI1.XI5.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<14>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<13>.MM_i_0 VSS! XI0.XI1.XI5.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<13>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<13>.MM_i_0_15 VSS! REG_DATA_9<13> XI0.XI1.XI5.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<13>.MM_i_0_15_63 XI0.XI1.XI5.XI3<13>.DUMMY1 REG_DATA_9<13>
+ XI0.XI1.XI5.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<13>.NEN
+ XI0.XI1.XI5.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<13>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<13>.MM_i_24 VDD! XI0.XI1.XI5.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<13>.MM_i_24_1 XI0.XI1.XI5.XI3<13>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<13>.MM_i_24_0 VDD! REG_DATA_9<13> XI0.XI1.XI5.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI5.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_9<13> XI0.XI1.XI5.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<13>.MM_i_24_1_48 XI0.XI1.XI5.XI3<13>.Y XI0.XI1.XI5.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<13>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI5.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI5.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI5.XI3<12>.MM_i_0 VSS! XI0.XI1.XI5.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI5.XI3<12>.MM_i_0_14 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<12>.MM_i_0_15 VSS! REG_DATA_9<12> XI0.XI1.XI5.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<12>.MM_i_0_15_63 XI0.XI1.XI5.XI3<12>.DUMMY1 REG_DATA_9<12>
+ XI0.XI1.XI5.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI5.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI5.XI3<12>.NEN
+ XI0.XI1.XI5.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI5.XI3<12>.MM_i_17 VSS! XI0.NET1<3> XI0.XI1.XI5.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI5.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI5.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<12>.MM_i_24 VDD! XI0.XI1.XI5.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI5.XI3<12>.MM_i_24_1 XI0.XI1.XI5.XI3<12>.DUMMY0 XI0.NET1<3>
+ XI0.XI1.XI5.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI5.XI3<12>.MM_i_24_0 VDD! REG_DATA_9<12> XI0.XI1.XI5.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI5.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_9<12> XI0.XI1.XI5.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI5.XI3<12>.MM_i_24_1_48 XI0.XI1.XI5.XI3<12>.Y XI0.XI1.XI5.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI5.XI3<12>.MM_i_42 VDD! XI0.NET1<3> XI0.XI1.XI5.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<3>.MM_i_0 VSS! XI0.XI1.XI10.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<3>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<3>.MM_i_0_15 VSS! REG_DATA_8<3> XI0.XI1.XI10.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<3>.MM_i_0_15_63 XI0.XI1.XI10.XI3<3>.DUMMY1 REG_DATA_8<3>
+ XI0.XI1.XI10.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<3>.NEN
+ XI0.XI1.XI10.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<3>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<3>.MM_i_24 VDD! XI0.XI1.XI10.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<3>.MM_i_24_1 XI0.XI1.XI10.XI3<3>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<3>.MM_i_24_0 VDD! REG_DATA_8<3> XI0.XI1.XI10.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_8<3> XI0.XI1.XI10.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<3>.MM_i_24_1_48 XI0.XI1.XI10.XI3<3>.Y XI0.XI1.XI10.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<3>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<2>.MM_i_0 VSS! XI0.XI1.XI10.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<2>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<2>.MM_i_0_15 VSS! REG_DATA_8<2> XI0.XI1.XI10.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<2>.MM_i_0_15_63 XI0.XI1.XI10.XI3<2>.DUMMY1 REG_DATA_8<2>
+ XI0.XI1.XI10.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<2>.NEN
+ XI0.XI1.XI10.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<2>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<2>.MM_i_24 VDD! XI0.XI1.XI10.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<2>.MM_i_24_1 XI0.XI1.XI10.XI3<2>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<2>.MM_i_24_0 VDD! REG_DATA_8<2> XI0.XI1.XI10.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_8<2> XI0.XI1.XI10.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<2>.MM_i_24_1_48 XI0.XI1.XI10.XI3<2>.Y XI0.XI1.XI10.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<2>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<1>.MM_i_0 VSS! XI0.XI1.XI10.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<1>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<1>.MM_i_0_15 VSS! REG_DATA_8<1> XI0.XI1.XI10.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<1>.MM_i_0_15_63 XI0.XI1.XI10.XI3<1>.DUMMY1 REG_DATA_8<1>
+ XI0.XI1.XI10.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<1>.NEN
+ XI0.XI1.XI10.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<1>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<1>.MM_i_24 VDD! XI0.XI1.XI10.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<1>.MM_i_24_1 XI0.XI1.XI10.XI3<1>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<1>.MM_i_24_0 VDD! REG_DATA_8<1> XI0.XI1.XI10.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_8<1> XI0.XI1.XI10.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<1>.MM_i_24_1_48 XI0.XI1.XI10.XI3<1>.Y XI0.XI1.XI10.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<1>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<0>.MM_i_0 VSS! XI0.XI1.XI10.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<0>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<0>.MM_i_0_15 VSS! REG_DATA_8<0> XI0.XI1.XI10.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<0>.MM_i_0_15_63 XI0.XI1.XI10.XI3<0>.DUMMY1 REG_DATA_8<0>
+ XI0.XI1.XI10.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<0>.NEN
+ XI0.XI1.XI10.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<0>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<0>.MM_i_24 VDD! XI0.XI1.XI10.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<0>.MM_i_24_1 XI0.XI1.XI10.XI3<0>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<0>.MM_i_24_0 VDD! REG_DATA_8<0> XI0.XI1.XI10.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_8<0> XI0.XI1.XI10.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<0>.MM_i_24_1_48 XI0.XI1.XI10.XI3<0>.Y XI0.XI1.XI10.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<0>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<7>.MM_i_0 VSS! XI0.XI1.XI10.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<7>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<7>.MM_i_0_15 VSS! REG_DATA_8<7> XI0.XI1.XI10.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<7>.MM_i_0_15_63 XI0.XI1.XI10.XI3<7>.DUMMY1 REG_DATA_8<7>
+ XI0.XI1.XI10.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<7>.NEN
+ XI0.XI1.XI10.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<7>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<7>.MM_i_24 VDD! XI0.XI1.XI10.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<7>.MM_i_24_1 XI0.XI1.XI10.XI3<7>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<7>.MM_i_24_0 VDD! REG_DATA_8<7> XI0.XI1.XI10.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_8<7> XI0.XI1.XI10.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<7>.MM_i_24_1_48 XI0.XI1.XI10.XI3<7>.Y XI0.XI1.XI10.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<7>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<6>.MM_i_0 VSS! XI0.XI1.XI10.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<6>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<6>.MM_i_0_15 VSS! REG_DATA_8<6> XI0.XI1.XI10.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<6>.MM_i_0_15_63 XI0.XI1.XI10.XI3<6>.DUMMY1 REG_DATA_8<6>
+ XI0.XI1.XI10.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<6>.NEN
+ XI0.XI1.XI10.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<6>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<6>.MM_i_24 VDD! XI0.XI1.XI10.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<6>.MM_i_24_1 XI0.XI1.XI10.XI3<6>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<6>.MM_i_24_0 VDD! REG_DATA_8<6> XI0.XI1.XI10.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_8<6> XI0.XI1.XI10.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<6>.MM_i_24_1_48 XI0.XI1.XI10.XI3<6>.Y XI0.XI1.XI10.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<6>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<5>.MM_i_0 VSS! XI0.XI1.XI10.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<5>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<5>.MM_i_0_15 VSS! REG_DATA_8<5> XI0.XI1.XI10.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<5>.MM_i_0_15_63 XI0.XI1.XI10.XI3<5>.DUMMY1 REG_DATA_8<5>
+ XI0.XI1.XI10.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<5>.NEN
+ XI0.XI1.XI10.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<5>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<5>.MM_i_24 VDD! XI0.XI1.XI10.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<5>.MM_i_24_1 XI0.XI1.XI10.XI3<5>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<5>.MM_i_24_0 VDD! REG_DATA_8<5> XI0.XI1.XI10.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_8<5> XI0.XI1.XI10.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<5>.MM_i_24_1_48 XI0.XI1.XI10.XI3<5>.Y XI0.XI1.XI10.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<5>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<4>.MM_i_0 VSS! XI0.XI1.XI10.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<4>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<4>.MM_i_0_15 VSS! REG_DATA_8<4> XI0.XI1.XI10.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<4>.MM_i_0_15_63 XI0.XI1.XI10.XI3<4>.DUMMY1 REG_DATA_8<4>
+ XI0.XI1.XI10.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<4>.NEN
+ XI0.XI1.XI10.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<4>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<4>.MM_i_24 VDD! XI0.XI1.XI10.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<4>.MM_i_24_1 XI0.XI1.XI10.XI3<4>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<4>.MM_i_24_0 VDD! REG_DATA_8<4> XI0.XI1.XI10.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_8<4> XI0.XI1.XI10.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<4>.MM_i_24_1_48 XI0.XI1.XI10.XI3<4>.Y XI0.XI1.XI10.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<4>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<11>.MM_i_0 VSS! XI0.XI1.XI10.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<11>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<11>.MM_i_0_15 VSS! REG_DATA_8<11> XI0.XI1.XI10.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<11>.MM_i_0_15_63 XI0.XI1.XI10.XI3<11>.DUMMY1 REG_DATA_8<11>
+ XI0.XI1.XI10.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<11>.NEN
+ XI0.XI1.XI10.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<11>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<11>.MM_i_24 VDD! XI0.XI1.XI10.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<11>.MM_i_24_1 XI0.XI1.XI10.XI3<11>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<11>.MM_i_24_0 VDD! REG_DATA_8<11> XI0.XI1.XI10.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_8<11> XI0.XI1.XI10.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<11>.MM_i_24_1_48 XI0.XI1.XI10.XI3<11>.Y
+ XI0.XI1.XI10.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI10.XI3<11>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<10>.MM_i_0 VSS! XI0.XI1.XI10.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<10>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<10>.MM_i_0_15 VSS! REG_DATA_8<10> XI0.XI1.XI10.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<10>.MM_i_0_15_63 XI0.XI1.XI10.XI3<10>.DUMMY1 REG_DATA_8<10>
+ XI0.XI1.XI10.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<10>.NEN
+ XI0.XI1.XI10.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<10>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<10>.MM_i_24 VDD! XI0.XI1.XI10.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<10>.MM_i_24_1 XI0.XI1.XI10.XI3<10>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<10>.MM_i_24_0 VDD! REG_DATA_8<10> XI0.XI1.XI10.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_8<10> XI0.XI1.XI10.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<10>.MM_i_24_1_48 XI0.XI1.XI10.XI3<10>.Y
+ XI0.XI1.XI10.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI10.XI3<10>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<9>.MM_i_0 VSS! XI0.XI1.XI10.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<9>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<9>.MM_i_0_15 VSS! REG_DATA_8<9> XI0.XI1.XI10.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<9>.MM_i_0_15_63 XI0.XI1.XI10.XI3<9>.DUMMY1 REG_DATA_8<9>
+ XI0.XI1.XI10.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<9>.NEN
+ XI0.XI1.XI10.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<9>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<9>.MM_i_24 VDD! XI0.XI1.XI10.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<9>.MM_i_24_1 XI0.XI1.XI10.XI3<9>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<9>.MM_i_24_0 VDD! REG_DATA_8<9> XI0.XI1.XI10.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_8<9> XI0.XI1.XI10.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<9>.MM_i_24_1_48 XI0.XI1.XI10.XI3<9>.Y XI0.XI1.XI10.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<9>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<8>.MM_i_0 VSS! XI0.XI1.XI10.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<8>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<8>.MM_i_0_15 VSS! REG_DATA_8<8> XI0.XI1.XI10.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<8>.MM_i_0_15_63 XI0.XI1.XI10.XI3<8>.DUMMY1 REG_DATA_8<8>
+ XI0.XI1.XI10.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<8>.NEN
+ XI0.XI1.XI10.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<8>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<8>.MM_i_24 VDD! XI0.XI1.XI10.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<8>.MM_i_24_1 XI0.XI1.XI10.XI3<8>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<8>.MM_i_24_0 VDD! REG_DATA_8<8> XI0.XI1.XI10.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_8<8> XI0.XI1.XI10.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI10.XI3<8>.MM_i_24_1_48 XI0.XI1.XI10.XI3<8>.Y XI0.XI1.XI10.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI10.XI3<8>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<15>.MM_i_0 VSS! XI0.XI1.XI10.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<15>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<15>.MM_i_0_15 VSS! REG_DATA_8<15> XI0.XI1.XI10.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<15>.MM_i_0_15_63 XI0.XI1.XI10.XI3<15>.DUMMY1 REG_DATA_8<15>
+ XI0.XI1.XI10.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<15>.NEN
+ XI0.XI1.XI10.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<15>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<15>.MM_i_24 VDD! XI0.XI1.XI10.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<15>.MM_i_24_1 XI0.XI1.XI10.XI3<15>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<15>.MM_i_24_0 VDD! REG_DATA_8<15> XI0.XI1.XI10.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_8<15> XI0.XI1.XI10.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<15>.MM_i_24_1_48 XI0.XI1.XI10.XI3<15>.Y
+ XI0.XI1.XI10.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI10.XI3<15>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<14>.MM_i_0 VSS! XI0.XI1.XI10.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<14>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<14>.MM_i_0_15 VSS! REG_DATA_8<14> XI0.XI1.XI10.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<14>.MM_i_0_15_63 XI0.XI1.XI10.XI3<14>.DUMMY1 REG_DATA_8<14>
+ XI0.XI1.XI10.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<14>.NEN
+ XI0.XI1.XI10.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<14>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<14>.MM_i_24 VDD! XI0.XI1.XI10.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<14>.MM_i_24_1 XI0.XI1.XI10.XI3<14>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<14>.MM_i_24_0 VDD! REG_DATA_8<14> XI0.XI1.XI10.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_8<14> XI0.XI1.XI10.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<14>.MM_i_24_1_48 XI0.XI1.XI10.XI3<14>.Y
+ XI0.XI1.XI10.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI10.XI3<14>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<13>.MM_i_0 VSS! XI0.XI1.XI10.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<13>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<13>.MM_i_0_15 VSS! REG_DATA_8<13> XI0.XI1.XI10.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<13>.MM_i_0_15_63 XI0.XI1.XI10.XI3<13>.DUMMY1 REG_DATA_8<13>
+ XI0.XI1.XI10.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<13>.NEN
+ XI0.XI1.XI10.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<13>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<13>.MM_i_24 VDD! XI0.XI1.XI10.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<13>.MM_i_24_1 XI0.XI1.XI10.XI3<13>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<13>.MM_i_24_0 VDD! REG_DATA_8<13> XI0.XI1.XI10.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_8<13> XI0.XI1.XI10.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<13>.MM_i_24_1_48 XI0.XI1.XI10.XI3<13>.Y
+ XI0.XI1.XI10.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI10.XI3<13>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI10.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI10.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI10.XI3<12>.MM_i_0 VSS! XI0.XI1.XI10.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI10.XI3<12>.MM_i_0_14 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<12>.MM_i_0_15 VSS! REG_DATA_8<12> XI0.XI1.XI10.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<12>.MM_i_0_15_63 XI0.XI1.XI10.XI3<12>.DUMMY1 REG_DATA_8<12>
+ XI0.XI1.XI10.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI10.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI10.XI3<12>.NEN
+ XI0.XI1.XI10.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI10.XI3<12>.MM_i_17 VSS! XI0.NET1<4> XI0.XI1.XI10.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI10.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI10.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<12>.MM_i_24 VDD! XI0.XI1.XI10.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI10.XI3<12>.MM_i_24_1 XI0.XI1.XI10.XI3<12>.DUMMY0 XI0.NET1<4>
+ XI0.XI1.XI10.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI10.XI3<12>.MM_i_24_0 VDD! REG_DATA_8<12> XI0.XI1.XI10.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_8<12> XI0.XI1.XI10.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI10.XI3<12>.MM_i_24_1_48 XI0.XI1.XI10.XI3<12>.Y
+ XI0.XI1.XI10.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI10.XI3<12>.MM_i_42 VDD! XI0.NET1<4> XI0.XI1.XI10.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<3>.MM_i_0 VSS! XI0.XI1.XI9.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<3>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<3>.MM_i_0_15 VSS! REG_DATA_7<3> XI0.XI1.XI9.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<3>.MM_i_0_15_63 XI0.XI1.XI9.XI3<3>.DUMMY1 REG_DATA_7<3>
+ XI0.XI1.XI9.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<3>.NEN
+ XI0.XI1.XI9.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<3>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<3>.MM_i_24 VDD! XI0.XI1.XI9.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<3>.MM_i_24_1 XI0.XI1.XI9.XI3<3>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<3>.MM_i_24_0 VDD! REG_DATA_7<3> XI0.XI1.XI9.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_7<3> XI0.XI1.XI9.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<3>.MM_i_24_1_48 XI0.XI1.XI9.XI3<3>.Y XI0.XI1.XI9.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<3>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<2>.MM_i_0 VSS! XI0.XI1.XI9.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<2>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<2>.MM_i_0_15 VSS! REG_DATA_7<2> XI0.XI1.XI9.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<2>.MM_i_0_15_63 XI0.XI1.XI9.XI3<2>.DUMMY1 REG_DATA_7<2>
+ XI0.XI1.XI9.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<2>.NEN
+ XI0.XI1.XI9.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<2>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<2>.MM_i_24 VDD! XI0.XI1.XI9.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<2>.MM_i_24_1 XI0.XI1.XI9.XI3<2>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<2>.MM_i_24_0 VDD! REG_DATA_7<2> XI0.XI1.XI9.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_7<2> XI0.XI1.XI9.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<2>.MM_i_24_1_48 XI0.XI1.XI9.XI3<2>.Y XI0.XI1.XI9.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<2>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<1>.MM_i_0 VSS! XI0.XI1.XI9.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<1>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<1>.MM_i_0_15 VSS! REG_DATA_7<1> XI0.XI1.XI9.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<1>.MM_i_0_15_63 XI0.XI1.XI9.XI3<1>.DUMMY1 REG_DATA_7<1>
+ XI0.XI1.XI9.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<1>.NEN
+ XI0.XI1.XI9.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<1>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<1>.MM_i_24 VDD! XI0.XI1.XI9.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<1>.MM_i_24_1 XI0.XI1.XI9.XI3<1>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<1>.MM_i_24_0 VDD! REG_DATA_7<1> XI0.XI1.XI9.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_7<1> XI0.XI1.XI9.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<1>.MM_i_24_1_48 XI0.XI1.XI9.XI3<1>.Y XI0.XI1.XI9.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<1>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<0>.MM_i_0 VSS! XI0.XI1.XI9.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<0>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<0>.MM_i_0_15 VSS! REG_DATA_7<0> XI0.XI1.XI9.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<0>.MM_i_0_15_63 XI0.XI1.XI9.XI3<0>.DUMMY1 REG_DATA_7<0>
+ XI0.XI1.XI9.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<0>.NEN
+ XI0.XI1.XI9.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<0>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<0>.MM_i_24 VDD! XI0.XI1.XI9.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<0>.MM_i_24_1 XI0.XI1.XI9.XI3<0>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<0>.MM_i_24_0 VDD! REG_DATA_7<0> XI0.XI1.XI9.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_7<0> XI0.XI1.XI9.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<0>.MM_i_24_1_48 XI0.XI1.XI9.XI3<0>.Y XI0.XI1.XI9.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<0>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<7>.MM_i_0 VSS! XI0.XI1.XI9.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<7>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<7>.MM_i_0_15 VSS! REG_DATA_7<7> XI0.XI1.XI9.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<7>.MM_i_0_15_63 XI0.XI1.XI9.XI3<7>.DUMMY1 REG_DATA_7<7>
+ XI0.XI1.XI9.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<7>.NEN
+ XI0.XI1.XI9.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<7>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<7>.MM_i_24 VDD! XI0.XI1.XI9.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<7>.MM_i_24_1 XI0.XI1.XI9.XI3<7>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<7>.MM_i_24_0 VDD! REG_DATA_7<7> XI0.XI1.XI9.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_7<7> XI0.XI1.XI9.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<7>.MM_i_24_1_48 XI0.XI1.XI9.XI3<7>.Y XI0.XI1.XI9.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<7>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<6>.MM_i_0 VSS! XI0.XI1.XI9.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<6>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<6>.MM_i_0_15 VSS! REG_DATA_7<6> XI0.XI1.XI9.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<6>.MM_i_0_15_63 XI0.XI1.XI9.XI3<6>.DUMMY1 REG_DATA_7<6>
+ XI0.XI1.XI9.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<6>.NEN
+ XI0.XI1.XI9.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<6>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<6>.MM_i_24 VDD! XI0.XI1.XI9.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<6>.MM_i_24_1 XI0.XI1.XI9.XI3<6>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<6>.MM_i_24_0 VDD! REG_DATA_7<6> XI0.XI1.XI9.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_7<6> XI0.XI1.XI9.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<6>.MM_i_24_1_48 XI0.XI1.XI9.XI3<6>.Y XI0.XI1.XI9.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<6>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<5>.MM_i_0 VSS! XI0.XI1.XI9.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<5>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<5>.MM_i_0_15 VSS! REG_DATA_7<5> XI0.XI1.XI9.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<5>.MM_i_0_15_63 XI0.XI1.XI9.XI3<5>.DUMMY1 REG_DATA_7<5>
+ XI0.XI1.XI9.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<5>.NEN
+ XI0.XI1.XI9.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<5>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<5>.MM_i_24 VDD! XI0.XI1.XI9.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<5>.MM_i_24_1 XI0.XI1.XI9.XI3<5>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<5>.MM_i_24_0 VDD! REG_DATA_7<5> XI0.XI1.XI9.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_7<5> XI0.XI1.XI9.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<5>.MM_i_24_1_48 XI0.XI1.XI9.XI3<5>.Y XI0.XI1.XI9.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<5>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<4>.MM_i_0 VSS! XI0.XI1.XI9.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<4>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<4>.MM_i_0_15 VSS! REG_DATA_7<4> XI0.XI1.XI9.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<4>.MM_i_0_15_63 XI0.XI1.XI9.XI3<4>.DUMMY1 REG_DATA_7<4>
+ XI0.XI1.XI9.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<4>.NEN
+ XI0.XI1.XI9.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<4>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<4>.MM_i_24 VDD! XI0.XI1.XI9.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<4>.MM_i_24_1 XI0.XI1.XI9.XI3<4>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<4>.MM_i_24_0 VDD! REG_DATA_7<4> XI0.XI1.XI9.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_7<4> XI0.XI1.XI9.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<4>.MM_i_24_1_48 XI0.XI1.XI9.XI3<4>.Y XI0.XI1.XI9.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<4>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<11>.MM_i_0 VSS! XI0.XI1.XI9.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<11>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<11>.MM_i_0_15 VSS! REG_DATA_7<11> XI0.XI1.XI9.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<11>.MM_i_0_15_63 XI0.XI1.XI9.XI3<11>.DUMMY1 REG_DATA_7<11>
+ XI0.XI1.XI9.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<11>.NEN
+ XI0.XI1.XI9.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<11>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<11>.MM_i_24 VDD! XI0.XI1.XI9.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<11>.MM_i_24_1 XI0.XI1.XI9.XI3<11>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<11>.MM_i_24_0 VDD! REG_DATA_7<11> XI0.XI1.XI9.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI9.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_7<11> XI0.XI1.XI9.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<11>.MM_i_24_1_48 XI0.XI1.XI9.XI3<11>.Y XI0.XI1.XI9.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<11>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<10>.MM_i_0 VSS! XI0.XI1.XI9.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<10>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<10>.MM_i_0_15 VSS! REG_DATA_7<10> XI0.XI1.XI9.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<10>.MM_i_0_15_63 XI0.XI1.XI9.XI3<10>.DUMMY1 REG_DATA_7<10>
+ XI0.XI1.XI9.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<10>.NEN
+ XI0.XI1.XI9.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<10>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<10>.MM_i_24 VDD! XI0.XI1.XI9.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<10>.MM_i_24_1 XI0.XI1.XI9.XI3<10>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<10>.MM_i_24_0 VDD! REG_DATA_7<10> XI0.XI1.XI9.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI9.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_7<10> XI0.XI1.XI9.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<10>.MM_i_24_1_48 XI0.XI1.XI9.XI3<10>.Y XI0.XI1.XI9.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<10>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<9>.MM_i_0 VSS! XI0.XI1.XI9.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<9>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<9>.MM_i_0_15 VSS! REG_DATA_7<9> XI0.XI1.XI9.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<9>.MM_i_0_15_63 XI0.XI1.XI9.XI3<9>.DUMMY1 REG_DATA_7<9>
+ XI0.XI1.XI9.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<9>.NEN
+ XI0.XI1.XI9.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<9>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<9>.MM_i_24 VDD! XI0.XI1.XI9.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<9>.MM_i_24_1 XI0.XI1.XI9.XI3<9>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<9>.MM_i_24_0 VDD! REG_DATA_7<9> XI0.XI1.XI9.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_7<9> XI0.XI1.XI9.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<9>.MM_i_24_1_48 XI0.XI1.XI9.XI3<9>.Y XI0.XI1.XI9.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<9>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<8>.MM_i_0 VSS! XI0.XI1.XI9.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<8>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<8>.MM_i_0_15 VSS! REG_DATA_7<8> XI0.XI1.XI9.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<8>.MM_i_0_15_63 XI0.XI1.XI9.XI3<8>.DUMMY1 REG_DATA_7<8>
+ XI0.XI1.XI9.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<8>.NEN
+ XI0.XI1.XI9.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<8>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<8>.MM_i_24 VDD! XI0.XI1.XI9.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<8>.MM_i_24_1 XI0.XI1.XI9.XI3<8>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<8>.MM_i_24_0 VDD! REG_DATA_7<8> XI0.XI1.XI9.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_7<8> XI0.XI1.XI9.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<8>.MM_i_24_1_48 XI0.XI1.XI9.XI3<8>.Y XI0.XI1.XI9.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<8>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<15>.MM_i_0 VSS! XI0.XI1.XI9.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<15>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<15>.MM_i_0_15 VSS! REG_DATA_7<15> XI0.XI1.XI9.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<15>.MM_i_0_15_63 XI0.XI1.XI9.XI3<15>.DUMMY1 REG_DATA_7<15>
+ XI0.XI1.XI9.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<15>.NEN
+ XI0.XI1.XI9.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<15>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<15>.MM_i_24 VDD! XI0.XI1.XI9.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<15>.MM_i_24_1 XI0.XI1.XI9.XI3<15>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<15>.MM_i_24_0 VDD! REG_DATA_7<15> XI0.XI1.XI9.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI9.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_7<15> XI0.XI1.XI9.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<15>.MM_i_24_1_48 XI0.XI1.XI9.XI3<15>.Y XI0.XI1.XI9.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<15>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<14>.MM_i_0 VSS! XI0.XI1.XI9.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<14>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<14>.MM_i_0_15 VSS! REG_DATA_7<14> XI0.XI1.XI9.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<14>.MM_i_0_15_63 XI0.XI1.XI9.XI3<14>.DUMMY1 REG_DATA_7<14>
+ XI0.XI1.XI9.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<14>.NEN
+ XI0.XI1.XI9.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<14>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<14>.MM_i_24 VDD! XI0.XI1.XI9.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<14>.MM_i_24_1 XI0.XI1.XI9.XI3<14>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<14>.MM_i_24_0 VDD! REG_DATA_7<14> XI0.XI1.XI9.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI9.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_7<14> XI0.XI1.XI9.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<14>.MM_i_24_1_48 XI0.XI1.XI9.XI3<14>.Y XI0.XI1.XI9.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<14>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<13>.MM_i_0 VSS! XI0.XI1.XI9.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<13>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<13>.MM_i_0_15 VSS! REG_DATA_7<13> XI0.XI1.XI9.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<13>.MM_i_0_15_63 XI0.XI1.XI9.XI3<13>.DUMMY1 REG_DATA_7<13>
+ XI0.XI1.XI9.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<13>.NEN
+ XI0.XI1.XI9.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<13>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<13>.MM_i_24 VDD! XI0.XI1.XI9.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<13>.MM_i_24_1 XI0.XI1.XI9.XI3<13>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<13>.MM_i_24_0 VDD! REG_DATA_7<13> XI0.XI1.XI9.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI9.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_7<13> XI0.XI1.XI9.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<13>.MM_i_24_1_48 XI0.XI1.XI9.XI3<13>.Y XI0.XI1.XI9.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<13>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI9.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI9.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI9.XI3<12>.MM_i_0 VSS! XI0.XI1.XI9.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI9.XI3<12>.MM_i_0_14 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<12>.MM_i_0_15 VSS! REG_DATA_7<12> XI0.XI1.XI9.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<12>.MM_i_0_15_63 XI0.XI1.XI9.XI3<12>.DUMMY1 REG_DATA_7<12>
+ XI0.XI1.XI9.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI9.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI9.XI3<12>.NEN
+ XI0.XI1.XI9.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI9.XI3<12>.MM_i_17 VSS! XI0.NET1<5> XI0.XI1.XI9.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI9.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI9.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<12>.MM_i_24 VDD! XI0.XI1.XI9.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI9.XI3<12>.MM_i_24_1 XI0.XI1.XI9.XI3<12>.DUMMY0 XI0.NET1<5>
+ XI0.XI1.XI9.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI9.XI3<12>.MM_i_24_0 VDD! REG_DATA_7<12> XI0.XI1.XI9.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI9.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_7<12> XI0.XI1.XI9.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI9.XI3<12>.MM_i_24_1_48 XI0.XI1.XI9.XI3<12>.Y XI0.XI1.XI9.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI9.XI3<12>.MM_i_42 VDD! XI0.NET1<5> XI0.XI1.XI9.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<3>.MM_i_0 VSS! XI0.XI1.XI7.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<3>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<3>.MM_i_0_15 VSS! REG_DATA_6<3> XI0.XI1.XI7.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<3>.MM_i_0_15_63 XI0.XI1.XI7.XI3<3>.DUMMY1 REG_DATA_6<3>
+ XI0.XI1.XI7.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<3>.NEN
+ XI0.XI1.XI7.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<3>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<3>.MM_i_24 VDD! XI0.XI1.XI7.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<3>.MM_i_24_1 XI0.XI1.XI7.XI3<3>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<3>.MM_i_24_0 VDD! REG_DATA_6<3> XI0.XI1.XI7.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_6<3> XI0.XI1.XI7.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<3>.MM_i_24_1_48 XI0.XI1.XI7.XI3<3>.Y XI0.XI1.XI7.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<3>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<2>.MM_i_0 VSS! XI0.XI1.XI7.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<2>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<2>.MM_i_0_15 VSS! REG_DATA_6<2> XI0.XI1.XI7.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<2>.MM_i_0_15_63 XI0.XI1.XI7.XI3<2>.DUMMY1 REG_DATA_6<2>
+ XI0.XI1.XI7.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<2>.NEN
+ XI0.XI1.XI7.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<2>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<2>.MM_i_24 VDD! XI0.XI1.XI7.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<2>.MM_i_24_1 XI0.XI1.XI7.XI3<2>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<2>.MM_i_24_0 VDD! REG_DATA_6<2> XI0.XI1.XI7.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_6<2> XI0.XI1.XI7.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<2>.MM_i_24_1_48 XI0.XI1.XI7.XI3<2>.Y XI0.XI1.XI7.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<2>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<1>.MM_i_0 VSS! XI0.XI1.XI7.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<1>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<1>.MM_i_0_15 VSS! REG_DATA_6<1> XI0.XI1.XI7.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<1>.MM_i_0_15_63 XI0.XI1.XI7.XI3<1>.DUMMY1 REG_DATA_6<1>
+ XI0.XI1.XI7.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<1>.NEN
+ XI0.XI1.XI7.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<1>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<1>.MM_i_24 VDD! XI0.XI1.XI7.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<1>.MM_i_24_1 XI0.XI1.XI7.XI3<1>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<1>.MM_i_24_0 VDD! REG_DATA_6<1> XI0.XI1.XI7.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_6<1> XI0.XI1.XI7.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<1>.MM_i_24_1_48 XI0.XI1.XI7.XI3<1>.Y XI0.XI1.XI7.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<1>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<0>.MM_i_0 VSS! XI0.XI1.XI7.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<0>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<0>.MM_i_0_15 VSS! REG_DATA_6<0> XI0.XI1.XI7.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<0>.MM_i_0_15_63 XI0.XI1.XI7.XI3<0>.DUMMY1 REG_DATA_6<0>
+ XI0.XI1.XI7.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<0>.NEN
+ XI0.XI1.XI7.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<0>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<0>.MM_i_24 VDD! XI0.XI1.XI7.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<0>.MM_i_24_1 XI0.XI1.XI7.XI3<0>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<0>.MM_i_24_0 VDD! REG_DATA_6<0> XI0.XI1.XI7.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_6<0> XI0.XI1.XI7.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<0>.MM_i_24_1_48 XI0.XI1.XI7.XI3<0>.Y XI0.XI1.XI7.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<0>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<7>.MM_i_0 VSS! XI0.XI1.XI7.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<7>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<7>.MM_i_0_15 VSS! REG_DATA_6<7> XI0.XI1.XI7.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<7>.MM_i_0_15_63 XI0.XI1.XI7.XI3<7>.DUMMY1 REG_DATA_6<7>
+ XI0.XI1.XI7.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<7>.NEN
+ XI0.XI1.XI7.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<7>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<7>.MM_i_24 VDD! XI0.XI1.XI7.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<7>.MM_i_24_1 XI0.XI1.XI7.XI3<7>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<7>.MM_i_24_0 VDD! REG_DATA_6<7> XI0.XI1.XI7.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_6<7> XI0.XI1.XI7.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<7>.MM_i_24_1_48 XI0.XI1.XI7.XI3<7>.Y XI0.XI1.XI7.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<7>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<6>.MM_i_0 VSS! XI0.XI1.XI7.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<6>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<6>.MM_i_0_15 VSS! REG_DATA_6<6> XI0.XI1.XI7.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<6>.MM_i_0_15_63 XI0.XI1.XI7.XI3<6>.DUMMY1 REG_DATA_6<6>
+ XI0.XI1.XI7.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<6>.NEN
+ XI0.XI1.XI7.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<6>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<6>.MM_i_24 VDD! XI0.XI1.XI7.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<6>.MM_i_24_1 XI0.XI1.XI7.XI3<6>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<6>.MM_i_24_0 VDD! REG_DATA_6<6> XI0.XI1.XI7.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_6<6> XI0.XI1.XI7.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<6>.MM_i_24_1_48 XI0.XI1.XI7.XI3<6>.Y XI0.XI1.XI7.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<6>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<5>.MM_i_0 VSS! XI0.XI1.XI7.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<5>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<5>.MM_i_0_15 VSS! REG_DATA_6<5> XI0.XI1.XI7.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<5>.MM_i_0_15_63 XI0.XI1.XI7.XI3<5>.DUMMY1 REG_DATA_6<5>
+ XI0.XI1.XI7.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<5>.NEN
+ XI0.XI1.XI7.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<5>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<5>.MM_i_24 VDD! XI0.XI1.XI7.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<5>.MM_i_24_1 XI0.XI1.XI7.XI3<5>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<5>.MM_i_24_0 VDD! REG_DATA_6<5> XI0.XI1.XI7.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_6<5> XI0.XI1.XI7.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<5>.MM_i_24_1_48 XI0.XI1.XI7.XI3<5>.Y XI0.XI1.XI7.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<5>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<4>.MM_i_0 VSS! XI0.XI1.XI7.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<4>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<4>.MM_i_0_15 VSS! REG_DATA_6<4> XI0.XI1.XI7.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<4>.MM_i_0_15_63 XI0.XI1.XI7.XI3<4>.DUMMY1 REG_DATA_6<4>
+ XI0.XI1.XI7.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<4>.NEN
+ XI0.XI1.XI7.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<4>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<4>.MM_i_24 VDD! XI0.XI1.XI7.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<4>.MM_i_24_1 XI0.XI1.XI7.XI3<4>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<4>.MM_i_24_0 VDD! REG_DATA_6<4> XI0.XI1.XI7.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_6<4> XI0.XI1.XI7.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<4>.MM_i_24_1_48 XI0.XI1.XI7.XI3<4>.Y XI0.XI1.XI7.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<4>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<11>.MM_i_0 VSS! XI0.XI1.XI7.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<11>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<11>.MM_i_0_15 VSS! REG_DATA_6<11> XI0.XI1.XI7.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<11>.MM_i_0_15_63 XI0.XI1.XI7.XI3<11>.DUMMY1 REG_DATA_6<11>
+ XI0.XI1.XI7.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<11>.NEN
+ XI0.XI1.XI7.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<11>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<11>.MM_i_24 VDD! XI0.XI1.XI7.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<11>.MM_i_24_1 XI0.XI1.XI7.XI3<11>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<11>.MM_i_24_0 VDD! REG_DATA_6<11> XI0.XI1.XI7.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI7.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_6<11> XI0.XI1.XI7.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<11>.MM_i_24_1_48 XI0.XI1.XI7.XI3<11>.Y XI0.XI1.XI7.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<11>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<10>.MM_i_0 VSS! XI0.XI1.XI7.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<10>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<10>.MM_i_0_15 VSS! REG_DATA_6<10> XI0.XI1.XI7.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<10>.MM_i_0_15_63 XI0.XI1.XI7.XI3<10>.DUMMY1 REG_DATA_6<10>
+ XI0.XI1.XI7.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<10>.NEN
+ XI0.XI1.XI7.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<10>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<10>.MM_i_24 VDD! XI0.XI1.XI7.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<10>.MM_i_24_1 XI0.XI1.XI7.XI3<10>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<10>.MM_i_24_0 VDD! REG_DATA_6<10> XI0.XI1.XI7.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI7.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_6<10> XI0.XI1.XI7.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<10>.MM_i_24_1_48 XI0.XI1.XI7.XI3<10>.Y XI0.XI1.XI7.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<10>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<9>.MM_i_0 VSS! XI0.XI1.XI7.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<9>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<9>.MM_i_0_15 VSS! REG_DATA_6<9> XI0.XI1.XI7.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<9>.MM_i_0_15_63 XI0.XI1.XI7.XI3<9>.DUMMY1 REG_DATA_6<9>
+ XI0.XI1.XI7.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<9>.NEN
+ XI0.XI1.XI7.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<9>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<9>.MM_i_24 VDD! XI0.XI1.XI7.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<9>.MM_i_24_1 XI0.XI1.XI7.XI3<9>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<9>.MM_i_24_0 VDD! REG_DATA_6<9> XI0.XI1.XI7.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_6<9> XI0.XI1.XI7.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<9>.MM_i_24_1_48 XI0.XI1.XI7.XI3<9>.Y XI0.XI1.XI7.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<9>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<8>.MM_i_0 VSS! XI0.XI1.XI7.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<8>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<8>.MM_i_0_15 VSS! REG_DATA_6<8> XI0.XI1.XI7.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<8>.MM_i_0_15_63 XI0.XI1.XI7.XI3<8>.DUMMY1 REG_DATA_6<8>
+ XI0.XI1.XI7.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<8>.NEN
+ XI0.XI1.XI7.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<8>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<8>.MM_i_24 VDD! XI0.XI1.XI7.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<8>.MM_i_24_1 XI0.XI1.XI7.XI3<8>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<8>.MM_i_24_0 VDD! REG_DATA_6<8> XI0.XI1.XI7.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_6<8> XI0.XI1.XI7.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<8>.MM_i_24_1_48 XI0.XI1.XI7.XI3<8>.Y XI0.XI1.XI7.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<8>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<15>.MM_i_0 VSS! XI0.XI1.XI7.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<15>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<15>.MM_i_0_15 VSS! REG_DATA_6<15> XI0.XI1.XI7.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<15>.MM_i_0_15_63 XI0.XI1.XI7.XI3<15>.DUMMY1 REG_DATA_6<15>
+ XI0.XI1.XI7.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<15>.NEN
+ XI0.XI1.XI7.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<15>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<15>.MM_i_24 VDD! XI0.XI1.XI7.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<15>.MM_i_24_1 XI0.XI1.XI7.XI3<15>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<15>.MM_i_24_0 VDD! REG_DATA_6<15> XI0.XI1.XI7.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI7.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_6<15> XI0.XI1.XI7.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<15>.MM_i_24_1_48 XI0.XI1.XI7.XI3<15>.Y XI0.XI1.XI7.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<15>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<14>.MM_i_0 VSS! XI0.XI1.XI7.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<14>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<14>.MM_i_0_15 VSS! REG_DATA_6<14> XI0.XI1.XI7.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<14>.MM_i_0_15_63 XI0.XI1.XI7.XI3<14>.DUMMY1 REG_DATA_6<14>
+ XI0.XI1.XI7.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<14>.NEN
+ XI0.XI1.XI7.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<14>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<14>.MM_i_24 VDD! XI0.XI1.XI7.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<14>.MM_i_24_1 XI0.XI1.XI7.XI3<14>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<14>.MM_i_24_0 VDD! REG_DATA_6<14> XI0.XI1.XI7.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI7.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_6<14> XI0.XI1.XI7.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<14>.MM_i_24_1_48 XI0.XI1.XI7.XI3<14>.Y XI0.XI1.XI7.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<14>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<13>.MM_i_0 VSS! XI0.XI1.XI7.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<13>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<13>.MM_i_0_15 VSS! REG_DATA_6<13> XI0.XI1.XI7.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<13>.MM_i_0_15_63 XI0.XI1.XI7.XI3<13>.DUMMY1 REG_DATA_6<13>
+ XI0.XI1.XI7.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<13>.NEN
+ XI0.XI1.XI7.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<13>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<13>.MM_i_24 VDD! XI0.XI1.XI7.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<13>.MM_i_24_1 XI0.XI1.XI7.XI3<13>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<13>.MM_i_24_0 VDD! REG_DATA_6<13> XI0.XI1.XI7.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI7.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_6<13> XI0.XI1.XI7.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<13>.MM_i_24_1_48 XI0.XI1.XI7.XI3<13>.Y XI0.XI1.XI7.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<13>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI7.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI7.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI7.XI3<12>.MM_i_0 VSS! XI0.XI1.XI7.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI7.XI3<12>.MM_i_0_14 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<12>.MM_i_0_15 VSS! REG_DATA_6<12> XI0.XI1.XI7.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<12>.MM_i_0_15_63 XI0.XI1.XI7.XI3<12>.DUMMY1 REG_DATA_6<12>
+ XI0.XI1.XI7.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI7.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI7.XI3<12>.NEN
+ XI0.XI1.XI7.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI7.XI3<12>.MM_i_17 VSS! XI0.NET1<6> XI0.XI1.XI7.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI7.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI7.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<12>.MM_i_24 VDD! XI0.XI1.XI7.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI7.XI3<12>.MM_i_24_1 XI0.XI1.XI7.XI3<12>.DUMMY0 XI0.NET1<6>
+ XI0.XI1.XI7.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI7.XI3<12>.MM_i_24_0 VDD! REG_DATA_6<12> XI0.XI1.XI7.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI7.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_6<12> XI0.XI1.XI7.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI7.XI3<12>.MM_i_24_1_48 XI0.XI1.XI7.XI3<12>.Y XI0.XI1.XI7.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI7.XI3<12>.MM_i_42 VDD! XI0.NET1<6> XI0.XI1.XI7.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<3>.MM_i_0 VSS! XI0.XI1.XI8.XI3<3>.X RD_DATA_0<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<3>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<3>.MM_i_0_15 VSS! REG_DATA_5<3> XI0.XI1.XI8.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<3>.MM_i_0_15_63 XI0.XI1.XI8.XI3<3>.DUMMY1 REG_DATA_5<3>
+ XI0.XI1.XI8.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<3>.NEN
+ XI0.XI1.XI8.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<3>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<3>.MM_i_24 VDD! XI0.XI1.XI8.XI3<3>.Y RD_DATA_0<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<3>.MM_i_24_1 XI0.XI1.XI8.XI3<3>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<3>.MM_i_24_0 VDD! REG_DATA_5<3> XI0.XI1.XI8.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_5<3> XI0.XI1.XI8.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<3>.MM_i_24_1_48 XI0.XI1.XI8.XI3<3>.Y XI0.XI1.XI8.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<3>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<2>.MM_i_0 VSS! XI0.XI1.XI8.XI3<2>.X RD_DATA_0<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<2>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<2>.MM_i_0_15 VSS! REG_DATA_5<2> XI0.XI1.XI8.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<2>.MM_i_0_15_63 XI0.XI1.XI8.XI3<2>.DUMMY1 REG_DATA_5<2>
+ XI0.XI1.XI8.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<2>.NEN
+ XI0.XI1.XI8.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<2>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<2>.MM_i_24 VDD! XI0.XI1.XI8.XI3<2>.Y RD_DATA_0<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<2>.MM_i_24_1 XI0.XI1.XI8.XI3<2>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<2>.MM_i_24_0 VDD! REG_DATA_5<2> XI0.XI1.XI8.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_5<2> XI0.XI1.XI8.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<2>.MM_i_24_1_48 XI0.XI1.XI8.XI3<2>.Y XI0.XI1.XI8.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<2>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<1>.MM_i_0 VSS! XI0.XI1.XI8.XI3<1>.X RD_DATA_0<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<1>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<1>.MM_i_0_15 VSS! REG_DATA_5<1> XI0.XI1.XI8.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<1>.MM_i_0_15_63 XI0.XI1.XI8.XI3<1>.DUMMY1 REG_DATA_5<1>
+ XI0.XI1.XI8.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<1>.NEN
+ XI0.XI1.XI8.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<1>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<1>.MM_i_24 VDD! XI0.XI1.XI8.XI3<1>.Y RD_DATA_0<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<1>.MM_i_24_1 XI0.XI1.XI8.XI3<1>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<1>.MM_i_24_0 VDD! REG_DATA_5<1> XI0.XI1.XI8.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_5<1> XI0.XI1.XI8.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<1>.MM_i_24_1_48 XI0.XI1.XI8.XI3<1>.Y XI0.XI1.XI8.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<1>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<0>.MM_i_0 VSS! XI0.XI1.XI8.XI3<0>.X RD_DATA_0<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<0>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<0>.MM_i_0_15 VSS! REG_DATA_5<0> XI0.XI1.XI8.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<0>.MM_i_0_15_63 XI0.XI1.XI8.XI3<0>.DUMMY1 REG_DATA_5<0>
+ XI0.XI1.XI8.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<0>.NEN
+ XI0.XI1.XI8.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<0>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<0>.MM_i_24 VDD! XI0.XI1.XI8.XI3<0>.Y RD_DATA_0<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<0>.MM_i_24_1 XI0.XI1.XI8.XI3<0>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<0>.MM_i_24_0 VDD! REG_DATA_5<0> XI0.XI1.XI8.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_5<0> XI0.XI1.XI8.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<0>.MM_i_24_1_48 XI0.XI1.XI8.XI3<0>.Y XI0.XI1.XI8.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<0>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<7>.MM_i_0 VSS! XI0.XI1.XI8.XI3<7>.X RD_DATA_0<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<7>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<7>.MM_i_0_15 VSS! REG_DATA_5<7> XI0.XI1.XI8.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<7>.MM_i_0_15_63 XI0.XI1.XI8.XI3<7>.DUMMY1 REG_DATA_5<7>
+ XI0.XI1.XI8.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<7>.NEN
+ XI0.XI1.XI8.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<7>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<7>.MM_i_24 VDD! XI0.XI1.XI8.XI3<7>.Y RD_DATA_0<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<7>.MM_i_24_1 XI0.XI1.XI8.XI3<7>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<7>.MM_i_24_0 VDD! REG_DATA_5<7> XI0.XI1.XI8.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_5<7> XI0.XI1.XI8.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<7>.MM_i_24_1_48 XI0.XI1.XI8.XI3<7>.Y XI0.XI1.XI8.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<7>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<6>.MM_i_0 VSS! XI0.XI1.XI8.XI3<6>.X RD_DATA_0<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<6>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<6>.MM_i_0_15 VSS! REG_DATA_5<6> XI0.XI1.XI8.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<6>.MM_i_0_15_63 XI0.XI1.XI8.XI3<6>.DUMMY1 REG_DATA_5<6>
+ XI0.XI1.XI8.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<6>.NEN
+ XI0.XI1.XI8.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<6>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<6>.MM_i_24 VDD! XI0.XI1.XI8.XI3<6>.Y RD_DATA_0<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<6>.MM_i_24_1 XI0.XI1.XI8.XI3<6>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<6>.MM_i_24_0 VDD! REG_DATA_5<6> XI0.XI1.XI8.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_5<6> XI0.XI1.XI8.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<6>.MM_i_24_1_48 XI0.XI1.XI8.XI3<6>.Y XI0.XI1.XI8.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<6>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<5>.MM_i_0 VSS! XI0.XI1.XI8.XI3<5>.X RD_DATA_0<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<5>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<5>.MM_i_0_15 VSS! REG_DATA_5<5> XI0.XI1.XI8.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<5>.MM_i_0_15_63 XI0.XI1.XI8.XI3<5>.DUMMY1 REG_DATA_5<5>
+ XI0.XI1.XI8.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<5>.NEN
+ XI0.XI1.XI8.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<5>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<5>.MM_i_24 VDD! XI0.XI1.XI8.XI3<5>.Y RD_DATA_0<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<5>.MM_i_24_1 XI0.XI1.XI8.XI3<5>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<5>.MM_i_24_0 VDD! REG_DATA_5<5> XI0.XI1.XI8.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_5<5> XI0.XI1.XI8.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<5>.MM_i_24_1_48 XI0.XI1.XI8.XI3<5>.Y XI0.XI1.XI8.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<5>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<4>.MM_i_0 VSS! XI0.XI1.XI8.XI3<4>.X RD_DATA_0<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<4>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<4>.MM_i_0_15 VSS! REG_DATA_5<4> XI0.XI1.XI8.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<4>.MM_i_0_15_63 XI0.XI1.XI8.XI3<4>.DUMMY1 REG_DATA_5<4>
+ XI0.XI1.XI8.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<4>.NEN
+ XI0.XI1.XI8.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<4>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<4>.MM_i_24 VDD! XI0.XI1.XI8.XI3<4>.Y RD_DATA_0<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<4>.MM_i_24_1 XI0.XI1.XI8.XI3<4>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<4>.MM_i_24_0 VDD! REG_DATA_5<4> XI0.XI1.XI8.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_5<4> XI0.XI1.XI8.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<4>.MM_i_24_1_48 XI0.XI1.XI8.XI3<4>.Y XI0.XI1.XI8.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<4>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<11>.MM_i_0 VSS! XI0.XI1.XI8.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<11>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<11>.MM_i_0_15 VSS! REG_DATA_5<11> XI0.XI1.XI8.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<11>.MM_i_0_15_63 XI0.XI1.XI8.XI3<11>.DUMMY1 REG_DATA_5<11>
+ XI0.XI1.XI8.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<11>.NEN
+ XI0.XI1.XI8.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<11>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<11>.MM_i_24 VDD! XI0.XI1.XI8.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<11>.MM_i_24_1 XI0.XI1.XI8.XI3<11>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<11>.MM_i_24_0 VDD! REG_DATA_5<11> XI0.XI1.XI8.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI8.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_5<11> XI0.XI1.XI8.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<11>.MM_i_24_1_48 XI0.XI1.XI8.XI3<11>.Y XI0.XI1.XI8.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<11>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<10>.MM_i_0 VSS! XI0.XI1.XI8.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<10>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<10>.MM_i_0_15 VSS! REG_DATA_5<10> XI0.XI1.XI8.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<10>.MM_i_0_15_63 XI0.XI1.XI8.XI3<10>.DUMMY1 REG_DATA_5<10>
+ XI0.XI1.XI8.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<10>.NEN
+ XI0.XI1.XI8.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<10>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<10>.MM_i_24 VDD! XI0.XI1.XI8.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<10>.MM_i_24_1 XI0.XI1.XI8.XI3<10>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<10>.MM_i_24_0 VDD! REG_DATA_5<10> XI0.XI1.XI8.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI8.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_5<10> XI0.XI1.XI8.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<10>.MM_i_24_1_48 XI0.XI1.XI8.XI3<10>.Y XI0.XI1.XI8.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<10>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<9>.MM_i_0 VSS! XI0.XI1.XI8.XI3<9>.X RD_DATA_0<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<9>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<9>.MM_i_0_15 VSS! REG_DATA_5<9> XI0.XI1.XI8.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<9>.MM_i_0_15_63 XI0.XI1.XI8.XI3<9>.DUMMY1 REG_DATA_5<9>
+ XI0.XI1.XI8.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<9>.NEN
+ XI0.XI1.XI8.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<9>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<9>.MM_i_24 VDD! XI0.XI1.XI8.XI3<9>.Y RD_DATA_0<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<9>.MM_i_24_1 XI0.XI1.XI8.XI3<9>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<9>.MM_i_24_0 VDD! REG_DATA_5<9> XI0.XI1.XI8.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_5<9> XI0.XI1.XI8.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<9>.MM_i_24_1_48 XI0.XI1.XI8.XI3<9>.Y XI0.XI1.XI8.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<9>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<8>.MM_i_0 VSS! XI0.XI1.XI8.XI3<8>.X RD_DATA_0<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<8>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<8>.MM_i_0_15 VSS! REG_DATA_5<8> XI0.XI1.XI8.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<8>.MM_i_0_15_63 XI0.XI1.XI8.XI3<8>.DUMMY1 REG_DATA_5<8>
+ XI0.XI1.XI8.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<8>.NEN
+ XI0.XI1.XI8.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<8>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<8>.MM_i_24 VDD! XI0.XI1.XI8.XI3<8>.Y RD_DATA_0<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<8>.MM_i_24_1 XI0.XI1.XI8.XI3<8>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<8>.MM_i_24_0 VDD! REG_DATA_5<8> XI0.XI1.XI8.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_5<8> XI0.XI1.XI8.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<8>.MM_i_24_1_48 XI0.XI1.XI8.XI3<8>.Y XI0.XI1.XI8.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<8>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<15>.MM_i_0 VSS! XI0.XI1.XI8.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<15>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<15>.MM_i_0_15 VSS! REG_DATA_5<15> XI0.XI1.XI8.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<15>.MM_i_0_15_63 XI0.XI1.XI8.XI3<15>.DUMMY1 REG_DATA_5<15>
+ XI0.XI1.XI8.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<15>.NEN
+ XI0.XI1.XI8.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<15>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<15>.MM_i_24 VDD! XI0.XI1.XI8.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<15>.MM_i_24_1 XI0.XI1.XI8.XI3<15>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<15>.MM_i_24_0 VDD! REG_DATA_5<15> XI0.XI1.XI8.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI8.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_5<15> XI0.XI1.XI8.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<15>.MM_i_24_1_48 XI0.XI1.XI8.XI3<15>.Y XI0.XI1.XI8.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<15>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<14>.MM_i_0 VSS! XI0.XI1.XI8.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<14>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<14>.MM_i_0_15 VSS! REG_DATA_5<14> XI0.XI1.XI8.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<14>.MM_i_0_15_63 XI0.XI1.XI8.XI3<14>.DUMMY1 REG_DATA_5<14>
+ XI0.XI1.XI8.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<14>.NEN
+ XI0.XI1.XI8.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<14>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<14>.MM_i_24 VDD! XI0.XI1.XI8.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<14>.MM_i_24_1 XI0.XI1.XI8.XI3<14>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<14>.MM_i_24_0 VDD! REG_DATA_5<14> XI0.XI1.XI8.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI8.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_5<14> XI0.XI1.XI8.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<14>.MM_i_24_1_48 XI0.XI1.XI8.XI3<14>.Y XI0.XI1.XI8.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<14>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<13>.MM_i_0 VSS! XI0.XI1.XI8.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<13>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<13>.MM_i_0_15 VSS! REG_DATA_5<13> XI0.XI1.XI8.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<13>.MM_i_0_15_63 XI0.XI1.XI8.XI3<13>.DUMMY1 REG_DATA_5<13>
+ XI0.XI1.XI8.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<13>.NEN
+ XI0.XI1.XI8.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<13>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<13>.MM_i_24 VDD! XI0.XI1.XI8.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<13>.MM_i_24_1 XI0.XI1.XI8.XI3<13>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<13>.MM_i_24_0 VDD! REG_DATA_5<13> XI0.XI1.XI8.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI8.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_5<13> XI0.XI1.XI8.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<13>.MM_i_24_1_48 XI0.XI1.XI8.XI3<13>.Y XI0.XI1.XI8.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<13>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI8.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI8.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI8.XI3<12>.MM_i_0 VSS! XI0.XI1.XI8.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI8.XI3<12>.MM_i_0_14 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<12>.MM_i_0_15 VSS! REG_DATA_5<12> XI0.XI1.XI8.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<12>.MM_i_0_15_63 XI0.XI1.XI8.XI3<12>.DUMMY1 REG_DATA_5<12>
+ XI0.XI1.XI8.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI8.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI8.XI3<12>.NEN
+ XI0.XI1.XI8.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI8.XI3<12>.MM_i_17 VSS! XI0.NET1<7> XI0.XI1.XI8.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI8.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI8.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<12>.MM_i_24 VDD! XI0.XI1.XI8.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI8.XI3<12>.MM_i_24_1 XI0.XI1.XI8.XI3<12>.DUMMY0 XI0.NET1<7>
+ XI0.XI1.XI8.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI8.XI3<12>.MM_i_24_0 VDD! REG_DATA_5<12> XI0.XI1.XI8.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI8.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_5<12> XI0.XI1.XI8.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI8.XI3<12>.MM_i_24_1_48 XI0.XI1.XI8.XI3<12>.Y XI0.XI1.XI8.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI8.XI3<12>.MM_i_42 VDD! XI0.NET1<7> XI0.XI1.XI8.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<3>.MM_i_0 VSS! XI0.XI1.XI11.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<3>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<3>.MM_i_0_15 VSS! REG_DATA_4<3> XI0.XI1.XI11.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<3>.MM_i_0_15_63 XI0.XI1.XI11.XI3<3>.DUMMY1 REG_DATA_4<3>
+ XI0.XI1.XI11.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<3>.NEN
+ XI0.XI1.XI11.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<3>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<3>.MM_i_24 VDD! XI0.XI1.XI11.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<3>.MM_i_24_1 XI0.XI1.XI11.XI3<3>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<3>.MM_i_24_0 VDD! REG_DATA_4<3> XI0.XI1.XI11.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_4<3> XI0.XI1.XI11.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<3>.MM_i_24_1_48 XI0.XI1.XI11.XI3<3>.Y XI0.XI1.XI11.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<3>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<2>.MM_i_0 VSS! XI0.XI1.XI11.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<2>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<2>.MM_i_0_15 VSS! REG_DATA_4<2> XI0.XI1.XI11.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<2>.MM_i_0_15_63 XI0.XI1.XI11.XI3<2>.DUMMY1 REG_DATA_4<2>
+ XI0.XI1.XI11.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<2>.NEN
+ XI0.XI1.XI11.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<2>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<2>.MM_i_24 VDD! XI0.XI1.XI11.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<2>.MM_i_24_1 XI0.XI1.XI11.XI3<2>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<2>.MM_i_24_0 VDD! REG_DATA_4<2> XI0.XI1.XI11.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_4<2> XI0.XI1.XI11.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<2>.MM_i_24_1_48 XI0.XI1.XI11.XI3<2>.Y XI0.XI1.XI11.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<2>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<1>.MM_i_0 VSS! XI0.XI1.XI11.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<1>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<1>.MM_i_0_15 VSS! REG_DATA_4<1> XI0.XI1.XI11.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<1>.MM_i_0_15_63 XI0.XI1.XI11.XI3<1>.DUMMY1 REG_DATA_4<1>
+ XI0.XI1.XI11.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<1>.NEN
+ XI0.XI1.XI11.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<1>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<1>.MM_i_24 VDD! XI0.XI1.XI11.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<1>.MM_i_24_1 XI0.XI1.XI11.XI3<1>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<1>.MM_i_24_0 VDD! REG_DATA_4<1> XI0.XI1.XI11.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_4<1> XI0.XI1.XI11.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<1>.MM_i_24_1_48 XI0.XI1.XI11.XI3<1>.Y XI0.XI1.XI11.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<1>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<0>.MM_i_0 VSS! XI0.XI1.XI11.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<0>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<0>.MM_i_0_15 VSS! REG_DATA_4<0> XI0.XI1.XI11.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<0>.MM_i_0_15_63 XI0.XI1.XI11.XI3<0>.DUMMY1 REG_DATA_4<0>
+ XI0.XI1.XI11.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<0>.NEN
+ XI0.XI1.XI11.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<0>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<0>.MM_i_24 VDD! XI0.XI1.XI11.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<0>.MM_i_24_1 XI0.XI1.XI11.XI3<0>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<0>.MM_i_24_0 VDD! REG_DATA_4<0> XI0.XI1.XI11.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_4<0> XI0.XI1.XI11.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<0>.MM_i_24_1_48 XI0.XI1.XI11.XI3<0>.Y XI0.XI1.XI11.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<0>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<7>.MM_i_0 VSS! XI0.XI1.XI11.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<7>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<7>.MM_i_0_15 VSS! REG_DATA_4<7> XI0.XI1.XI11.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<7>.MM_i_0_15_63 XI0.XI1.XI11.XI3<7>.DUMMY1 REG_DATA_4<7>
+ XI0.XI1.XI11.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<7>.NEN
+ XI0.XI1.XI11.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<7>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<7>.MM_i_24 VDD! XI0.XI1.XI11.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<7>.MM_i_24_1 XI0.XI1.XI11.XI3<7>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<7>.MM_i_24_0 VDD! REG_DATA_4<7> XI0.XI1.XI11.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_4<7> XI0.XI1.XI11.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<7>.MM_i_24_1_48 XI0.XI1.XI11.XI3<7>.Y XI0.XI1.XI11.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<7>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<6>.MM_i_0 VSS! XI0.XI1.XI11.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<6>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<6>.MM_i_0_15 VSS! REG_DATA_4<6> XI0.XI1.XI11.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<6>.MM_i_0_15_63 XI0.XI1.XI11.XI3<6>.DUMMY1 REG_DATA_4<6>
+ XI0.XI1.XI11.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<6>.NEN
+ XI0.XI1.XI11.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<6>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<6>.MM_i_24 VDD! XI0.XI1.XI11.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<6>.MM_i_24_1 XI0.XI1.XI11.XI3<6>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<6>.MM_i_24_0 VDD! REG_DATA_4<6> XI0.XI1.XI11.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_4<6> XI0.XI1.XI11.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<6>.MM_i_24_1_48 XI0.XI1.XI11.XI3<6>.Y XI0.XI1.XI11.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<6>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<5>.MM_i_0 VSS! XI0.XI1.XI11.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<5>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<5>.MM_i_0_15 VSS! REG_DATA_4<5> XI0.XI1.XI11.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<5>.MM_i_0_15_63 XI0.XI1.XI11.XI3<5>.DUMMY1 REG_DATA_4<5>
+ XI0.XI1.XI11.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<5>.NEN
+ XI0.XI1.XI11.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<5>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<5>.MM_i_24 VDD! XI0.XI1.XI11.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<5>.MM_i_24_1 XI0.XI1.XI11.XI3<5>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<5>.MM_i_24_0 VDD! REG_DATA_4<5> XI0.XI1.XI11.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_4<5> XI0.XI1.XI11.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<5>.MM_i_24_1_48 XI0.XI1.XI11.XI3<5>.Y XI0.XI1.XI11.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<5>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<4>.MM_i_0 VSS! XI0.XI1.XI11.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<4>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<4>.MM_i_0_15 VSS! REG_DATA_4<4> XI0.XI1.XI11.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<4>.MM_i_0_15_63 XI0.XI1.XI11.XI3<4>.DUMMY1 REG_DATA_4<4>
+ XI0.XI1.XI11.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<4>.NEN
+ XI0.XI1.XI11.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<4>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<4>.MM_i_24 VDD! XI0.XI1.XI11.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<4>.MM_i_24_1 XI0.XI1.XI11.XI3<4>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<4>.MM_i_24_0 VDD! REG_DATA_4<4> XI0.XI1.XI11.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_4<4> XI0.XI1.XI11.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<4>.MM_i_24_1_48 XI0.XI1.XI11.XI3<4>.Y XI0.XI1.XI11.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<4>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<11>.MM_i_0 VSS! XI0.XI1.XI11.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<11>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<11>.MM_i_0_15 VSS! REG_DATA_4<11> XI0.XI1.XI11.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<11>.MM_i_0_15_63 XI0.XI1.XI11.XI3<11>.DUMMY1 REG_DATA_4<11>
+ XI0.XI1.XI11.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<11>.NEN
+ XI0.XI1.XI11.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<11>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<11>.MM_i_24 VDD! XI0.XI1.XI11.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<11>.MM_i_24_1 XI0.XI1.XI11.XI3<11>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<11>.MM_i_24_0 VDD! REG_DATA_4<11> XI0.XI1.XI11.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_4<11> XI0.XI1.XI11.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<11>.MM_i_24_1_48 XI0.XI1.XI11.XI3<11>.Y
+ XI0.XI1.XI11.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI11.XI3<11>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<10>.MM_i_0 VSS! XI0.XI1.XI11.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<10>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<10>.MM_i_0_15 VSS! REG_DATA_4<10> XI0.XI1.XI11.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<10>.MM_i_0_15_63 XI0.XI1.XI11.XI3<10>.DUMMY1 REG_DATA_4<10>
+ XI0.XI1.XI11.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<10>.NEN
+ XI0.XI1.XI11.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<10>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<10>.MM_i_24 VDD! XI0.XI1.XI11.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<10>.MM_i_24_1 XI0.XI1.XI11.XI3<10>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<10>.MM_i_24_0 VDD! REG_DATA_4<10> XI0.XI1.XI11.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_4<10> XI0.XI1.XI11.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<10>.MM_i_24_1_48 XI0.XI1.XI11.XI3<10>.Y
+ XI0.XI1.XI11.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI11.XI3<10>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<9>.MM_i_0 VSS! XI0.XI1.XI11.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<9>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<9>.MM_i_0_15 VSS! REG_DATA_4<9> XI0.XI1.XI11.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<9>.MM_i_0_15_63 XI0.XI1.XI11.XI3<9>.DUMMY1 REG_DATA_4<9>
+ XI0.XI1.XI11.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<9>.NEN
+ XI0.XI1.XI11.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<9>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<9>.MM_i_24 VDD! XI0.XI1.XI11.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<9>.MM_i_24_1 XI0.XI1.XI11.XI3<9>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<9>.MM_i_24_0 VDD! REG_DATA_4<9> XI0.XI1.XI11.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_4<9> XI0.XI1.XI11.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<9>.MM_i_24_1_48 XI0.XI1.XI11.XI3<9>.Y XI0.XI1.XI11.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<9>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<8>.MM_i_0 VSS! XI0.XI1.XI11.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<8>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<8>.MM_i_0_15 VSS! REG_DATA_4<8> XI0.XI1.XI11.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<8>.MM_i_0_15_63 XI0.XI1.XI11.XI3<8>.DUMMY1 REG_DATA_4<8>
+ XI0.XI1.XI11.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<8>.NEN
+ XI0.XI1.XI11.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<8>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<8>.MM_i_24 VDD! XI0.XI1.XI11.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<8>.MM_i_24_1 XI0.XI1.XI11.XI3<8>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<8>.MM_i_24_0 VDD! REG_DATA_4<8> XI0.XI1.XI11.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_4<8> XI0.XI1.XI11.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI11.XI3<8>.MM_i_24_1_48 XI0.XI1.XI11.XI3<8>.Y XI0.XI1.XI11.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI11.XI3<8>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<15>.MM_i_0 VSS! XI0.XI1.XI11.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<15>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<15>.MM_i_0_15 VSS! REG_DATA_4<15> XI0.XI1.XI11.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<15>.MM_i_0_15_63 XI0.XI1.XI11.XI3<15>.DUMMY1 REG_DATA_4<15>
+ XI0.XI1.XI11.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<15>.NEN
+ XI0.XI1.XI11.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<15>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<15>.MM_i_24 VDD! XI0.XI1.XI11.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<15>.MM_i_24_1 XI0.XI1.XI11.XI3<15>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<15>.MM_i_24_0 VDD! REG_DATA_4<15> XI0.XI1.XI11.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_4<15> XI0.XI1.XI11.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<15>.MM_i_24_1_48 XI0.XI1.XI11.XI3<15>.Y
+ XI0.XI1.XI11.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI11.XI3<15>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<14>.MM_i_0 VSS! XI0.XI1.XI11.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<14>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<14>.MM_i_0_15 VSS! REG_DATA_4<14> XI0.XI1.XI11.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<14>.MM_i_0_15_63 XI0.XI1.XI11.XI3<14>.DUMMY1 REG_DATA_4<14>
+ XI0.XI1.XI11.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<14>.NEN
+ XI0.XI1.XI11.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<14>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<14>.MM_i_24 VDD! XI0.XI1.XI11.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<14>.MM_i_24_1 XI0.XI1.XI11.XI3<14>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<14>.MM_i_24_0 VDD! REG_DATA_4<14> XI0.XI1.XI11.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_4<14> XI0.XI1.XI11.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<14>.MM_i_24_1_48 XI0.XI1.XI11.XI3<14>.Y
+ XI0.XI1.XI11.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI11.XI3<14>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<13>.MM_i_0 VSS! XI0.XI1.XI11.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<13>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<13>.MM_i_0_15 VSS! REG_DATA_4<13> XI0.XI1.XI11.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<13>.MM_i_0_15_63 XI0.XI1.XI11.XI3<13>.DUMMY1 REG_DATA_4<13>
+ XI0.XI1.XI11.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<13>.NEN
+ XI0.XI1.XI11.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<13>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<13>.MM_i_24 VDD! XI0.XI1.XI11.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<13>.MM_i_24_1 XI0.XI1.XI11.XI3<13>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<13>.MM_i_24_0 VDD! REG_DATA_4<13> XI0.XI1.XI11.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_4<13> XI0.XI1.XI11.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<13>.MM_i_24_1_48 XI0.XI1.XI11.XI3<13>.Y
+ XI0.XI1.XI11.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI11.XI3<13>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI11.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI11.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI11.XI3<12>.MM_i_0 VSS! XI0.XI1.XI11.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI11.XI3<12>.MM_i_0_14 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<12>.MM_i_0_15 VSS! REG_DATA_4<12> XI0.XI1.XI11.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<12>.MM_i_0_15_63 XI0.XI1.XI11.XI3<12>.DUMMY1 REG_DATA_4<12>
+ XI0.XI1.XI11.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI11.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI11.XI3<12>.NEN
+ XI0.XI1.XI11.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI11.XI3<12>.MM_i_17 VSS! XI0.NET1<8> XI0.XI1.XI11.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI11.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI11.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<12>.MM_i_24 VDD! XI0.XI1.XI11.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI11.XI3<12>.MM_i_24_1 XI0.XI1.XI11.XI3<12>.DUMMY0 XI0.NET1<8>
+ XI0.XI1.XI11.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI11.XI3<12>.MM_i_24_0 VDD! REG_DATA_4<12> XI0.XI1.XI11.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_4<12> XI0.XI1.XI11.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI11.XI3<12>.MM_i_24_1_48 XI0.XI1.XI11.XI3<12>.Y
+ XI0.XI1.XI11.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI11.XI3<12>.MM_i_42 VDD! XI0.NET1<8> XI0.XI1.XI11.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<3>.MM_i_0 VSS! XI0.XI1.XI12.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<3>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<3>.MM_i_0_15 VSS! REG_DATA_3<3> XI0.XI1.XI12.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<3>.MM_i_0_15_63 XI0.XI1.XI12.XI3<3>.DUMMY1 REG_DATA_3<3>
+ XI0.XI1.XI12.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<3>.NEN
+ XI0.XI1.XI12.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<3>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<3>.MM_i_24 VDD! XI0.XI1.XI12.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<3>.MM_i_24_1 XI0.XI1.XI12.XI3<3>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<3>.MM_i_24_0 VDD! REG_DATA_3<3> XI0.XI1.XI12.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_3<3> XI0.XI1.XI12.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<3>.MM_i_24_1_48 XI0.XI1.XI12.XI3<3>.Y XI0.XI1.XI12.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<3>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<2>.MM_i_0 VSS! XI0.XI1.XI12.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<2>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<2>.MM_i_0_15 VSS! REG_DATA_3<2> XI0.XI1.XI12.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<2>.MM_i_0_15_63 XI0.XI1.XI12.XI3<2>.DUMMY1 REG_DATA_3<2>
+ XI0.XI1.XI12.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<2>.NEN
+ XI0.XI1.XI12.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<2>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<2>.MM_i_24 VDD! XI0.XI1.XI12.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<2>.MM_i_24_1 XI0.XI1.XI12.XI3<2>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<2>.MM_i_24_0 VDD! REG_DATA_3<2> XI0.XI1.XI12.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_3<2> XI0.XI1.XI12.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<2>.MM_i_24_1_48 XI0.XI1.XI12.XI3<2>.Y XI0.XI1.XI12.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<2>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<1>.MM_i_0 VSS! XI0.XI1.XI12.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<1>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<1>.MM_i_0_15 VSS! REG_DATA_3<1> XI0.XI1.XI12.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<1>.MM_i_0_15_63 XI0.XI1.XI12.XI3<1>.DUMMY1 REG_DATA_3<1>
+ XI0.XI1.XI12.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<1>.NEN
+ XI0.XI1.XI12.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<1>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<1>.MM_i_24 VDD! XI0.XI1.XI12.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<1>.MM_i_24_1 XI0.XI1.XI12.XI3<1>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<1>.MM_i_24_0 VDD! REG_DATA_3<1> XI0.XI1.XI12.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_3<1> XI0.XI1.XI12.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<1>.MM_i_24_1_48 XI0.XI1.XI12.XI3<1>.Y XI0.XI1.XI12.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<1>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<0>.MM_i_0 VSS! XI0.XI1.XI12.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<0>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<0>.MM_i_0_15 VSS! REG_DATA_3<0> XI0.XI1.XI12.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<0>.MM_i_0_15_63 XI0.XI1.XI12.XI3<0>.DUMMY1 REG_DATA_3<0>
+ XI0.XI1.XI12.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<0>.NEN
+ XI0.XI1.XI12.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<0>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<0>.MM_i_24 VDD! XI0.XI1.XI12.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<0>.MM_i_24_1 XI0.XI1.XI12.XI3<0>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<0>.MM_i_24_0 VDD! REG_DATA_3<0> XI0.XI1.XI12.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_3<0> XI0.XI1.XI12.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<0>.MM_i_24_1_48 XI0.XI1.XI12.XI3<0>.Y XI0.XI1.XI12.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<0>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<7>.MM_i_0 VSS! XI0.XI1.XI12.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<7>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<7>.MM_i_0_15 VSS! REG_DATA_3<7> XI0.XI1.XI12.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<7>.MM_i_0_15_63 XI0.XI1.XI12.XI3<7>.DUMMY1 REG_DATA_3<7>
+ XI0.XI1.XI12.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<7>.NEN
+ XI0.XI1.XI12.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<7>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<7>.MM_i_24 VDD! XI0.XI1.XI12.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<7>.MM_i_24_1 XI0.XI1.XI12.XI3<7>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<7>.MM_i_24_0 VDD! REG_DATA_3<7> XI0.XI1.XI12.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_3<7> XI0.XI1.XI12.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<7>.MM_i_24_1_48 XI0.XI1.XI12.XI3<7>.Y XI0.XI1.XI12.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<7>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<6>.MM_i_0 VSS! XI0.XI1.XI12.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<6>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<6>.MM_i_0_15 VSS! REG_DATA_3<6> XI0.XI1.XI12.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<6>.MM_i_0_15_63 XI0.XI1.XI12.XI3<6>.DUMMY1 REG_DATA_3<6>
+ XI0.XI1.XI12.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<6>.NEN
+ XI0.XI1.XI12.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<6>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<6>.MM_i_24 VDD! XI0.XI1.XI12.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<6>.MM_i_24_1 XI0.XI1.XI12.XI3<6>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<6>.MM_i_24_0 VDD! REG_DATA_3<6> XI0.XI1.XI12.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_3<6> XI0.XI1.XI12.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<6>.MM_i_24_1_48 XI0.XI1.XI12.XI3<6>.Y XI0.XI1.XI12.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<6>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<5>.MM_i_0 VSS! XI0.XI1.XI12.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<5>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<5>.MM_i_0_15 VSS! REG_DATA_3<5> XI0.XI1.XI12.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<5>.MM_i_0_15_63 XI0.XI1.XI12.XI3<5>.DUMMY1 REG_DATA_3<5>
+ XI0.XI1.XI12.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<5>.NEN
+ XI0.XI1.XI12.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<5>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<5>.MM_i_24 VDD! XI0.XI1.XI12.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<5>.MM_i_24_1 XI0.XI1.XI12.XI3<5>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<5>.MM_i_24_0 VDD! REG_DATA_3<5> XI0.XI1.XI12.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_3<5> XI0.XI1.XI12.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<5>.MM_i_24_1_48 XI0.XI1.XI12.XI3<5>.Y XI0.XI1.XI12.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<5>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<4>.MM_i_0 VSS! XI0.XI1.XI12.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<4>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<4>.MM_i_0_15 VSS! REG_DATA_3<4> XI0.XI1.XI12.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<4>.MM_i_0_15_63 XI0.XI1.XI12.XI3<4>.DUMMY1 REG_DATA_3<4>
+ XI0.XI1.XI12.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<4>.NEN
+ XI0.XI1.XI12.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<4>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<4>.MM_i_24 VDD! XI0.XI1.XI12.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<4>.MM_i_24_1 XI0.XI1.XI12.XI3<4>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<4>.MM_i_24_0 VDD! REG_DATA_3<4> XI0.XI1.XI12.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_3<4> XI0.XI1.XI12.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<4>.MM_i_24_1_48 XI0.XI1.XI12.XI3<4>.Y XI0.XI1.XI12.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<4>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<11>.MM_i_0 VSS! XI0.XI1.XI12.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<11>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<11>.MM_i_0_15 VSS! REG_DATA_3<11> XI0.XI1.XI12.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<11>.MM_i_0_15_63 XI0.XI1.XI12.XI3<11>.DUMMY1 REG_DATA_3<11>
+ XI0.XI1.XI12.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<11>.NEN
+ XI0.XI1.XI12.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<11>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<11>.MM_i_24 VDD! XI0.XI1.XI12.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<11>.MM_i_24_1 XI0.XI1.XI12.XI3<11>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<11>.MM_i_24_0 VDD! REG_DATA_3<11> XI0.XI1.XI12.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_3<11> XI0.XI1.XI12.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<11>.MM_i_24_1_48 XI0.XI1.XI12.XI3<11>.Y
+ XI0.XI1.XI12.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI12.XI3<11>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<10>.MM_i_0 VSS! XI0.XI1.XI12.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<10>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<10>.MM_i_0_15 VSS! REG_DATA_3<10> XI0.XI1.XI12.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<10>.MM_i_0_15_63 XI0.XI1.XI12.XI3<10>.DUMMY1 REG_DATA_3<10>
+ XI0.XI1.XI12.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<10>.NEN
+ XI0.XI1.XI12.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<10>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<10>.MM_i_24 VDD! XI0.XI1.XI12.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<10>.MM_i_24_1 XI0.XI1.XI12.XI3<10>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<10>.MM_i_24_0 VDD! REG_DATA_3<10> XI0.XI1.XI12.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_3<10> XI0.XI1.XI12.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<10>.MM_i_24_1_48 XI0.XI1.XI12.XI3<10>.Y
+ XI0.XI1.XI12.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI12.XI3<10>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<9>.MM_i_0 VSS! XI0.XI1.XI12.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<9>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<9>.MM_i_0_15 VSS! REG_DATA_3<9> XI0.XI1.XI12.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<9>.MM_i_0_15_63 XI0.XI1.XI12.XI3<9>.DUMMY1 REG_DATA_3<9>
+ XI0.XI1.XI12.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<9>.NEN
+ XI0.XI1.XI12.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<9>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<9>.MM_i_24 VDD! XI0.XI1.XI12.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<9>.MM_i_24_1 XI0.XI1.XI12.XI3<9>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<9>.MM_i_24_0 VDD! REG_DATA_3<9> XI0.XI1.XI12.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_3<9> XI0.XI1.XI12.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<9>.MM_i_24_1_48 XI0.XI1.XI12.XI3<9>.Y XI0.XI1.XI12.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<9>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<8>.MM_i_0 VSS! XI0.XI1.XI12.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<8>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<8>.MM_i_0_15 VSS! REG_DATA_3<8> XI0.XI1.XI12.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<8>.MM_i_0_15_63 XI0.XI1.XI12.XI3<8>.DUMMY1 REG_DATA_3<8>
+ XI0.XI1.XI12.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<8>.NEN
+ XI0.XI1.XI12.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<8>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<8>.MM_i_24 VDD! XI0.XI1.XI12.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<8>.MM_i_24_1 XI0.XI1.XI12.XI3<8>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<8>.MM_i_24_0 VDD! REG_DATA_3<8> XI0.XI1.XI12.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_3<8> XI0.XI1.XI12.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI12.XI3<8>.MM_i_24_1_48 XI0.XI1.XI12.XI3<8>.Y XI0.XI1.XI12.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI12.XI3<8>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<15>.MM_i_0 VSS! XI0.XI1.XI12.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<15>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<15>.MM_i_0_15 VSS! REG_DATA_3<15> XI0.XI1.XI12.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<15>.MM_i_0_15_63 XI0.XI1.XI12.XI3<15>.DUMMY1 REG_DATA_3<15>
+ XI0.XI1.XI12.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<15>.NEN
+ XI0.XI1.XI12.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<15>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<15>.MM_i_24 VDD! XI0.XI1.XI12.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<15>.MM_i_24_1 XI0.XI1.XI12.XI3<15>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<15>.MM_i_24_0 VDD! REG_DATA_3<15> XI0.XI1.XI12.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_3<15> XI0.XI1.XI12.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<15>.MM_i_24_1_48 XI0.XI1.XI12.XI3<15>.Y
+ XI0.XI1.XI12.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI12.XI3<15>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<14>.MM_i_0 VSS! XI0.XI1.XI12.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<14>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<14>.MM_i_0_15 VSS! REG_DATA_3<14> XI0.XI1.XI12.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<14>.MM_i_0_15_63 XI0.XI1.XI12.XI3<14>.DUMMY1 REG_DATA_3<14>
+ XI0.XI1.XI12.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<14>.NEN
+ XI0.XI1.XI12.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<14>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<14>.MM_i_24 VDD! XI0.XI1.XI12.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<14>.MM_i_24_1 XI0.XI1.XI12.XI3<14>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<14>.MM_i_24_0 VDD! REG_DATA_3<14> XI0.XI1.XI12.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_3<14> XI0.XI1.XI12.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<14>.MM_i_24_1_48 XI0.XI1.XI12.XI3<14>.Y
+ XI0.XI1.XI12.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI12.XI3<14>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<13>.MM_i_0 VSS! XI0.XI1.XI12.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<13>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<13>.MM_i_0_15 VSS! REG_DATA_3<13> XI0.XI1.XI12.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<13>.MM_i_0_15_63 XI0.XI1.XI12.XI3<13>.DUMMY1 REG_DATA_3<13>
+ XI0.XI1.XI12.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<13>.NEN
+ XI0.XI1.XI12.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<13>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<13>.MM_i_24 VDD! XI0.XI1.XI12.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<13>.MM_i_24_1 XI0.XI1.XI12.XI3<13>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<13>.MM_i_24_0 VDD! REG_DATA_3<13> XI0.XI1.XI12.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_3<13> XI0.XI1.XI12.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<13>.MM_i_24_1_48 XI0.XI1.XI12.XI3<13>.Y
+ XI0.XI1.XI12.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI12.XI3<13>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI12.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI12.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI12.XI3<12>.MM_i_0 VSS! XI0.XI1.XI12.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI12.XI3<12>.MM_i_0_14 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<12>.MM_i_0_15 VSS! REG_DATA_3<12> XI0.XI1.XI12.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<12>.MM_i_0_15_63 XI0.XI1.XI12.XI3<12>.DUMMY1 REG_DATA_3<12>
+ XI0.XI1.XI12.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI12.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI12.XI3<12>.NEN
+ XI0.XI1.XI12.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI12.XI3<12>.MM_i_17 VSS! XI0.NET1<9> XI0.XI1.XI12.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI12.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI12.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<12>.MM_i_24 VDD! XI0.XI1.XI12.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI12.XI3<12>.MM_i_24_1 XI0.XI1.XI12.XI3<12>.DUMMY0 XI0.NET1<9>
+ XI0.XI1.XI12.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI12.XI3<12>.MM_i_24_0 VDD! REG_DATA_3<12> XI0.XI1.XI12.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_3<12> XI0.XI1.XI12.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI12.XI3<12>.MM_i_24_1_48 XI0.XI1.XI12.XI3<12>.Y
+ XI0.XI1.XI12.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI12.XI3<12>.MM_i_42 VDD! XI0.NET1<9> XI0.XI1.XI12.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<3>.MM_i_0 VSS! XI0.XI1.XI14.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<3>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<3>.MM_i_0_15 VSS! REG_DATA_2<3> XI0.XI1.XI14.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<3>.MM_i_0_15_63 XI0.XI1.XI14.XI3<3>.DUMMY1 REG_DATA_2<3>
+ XI0.XI1.XI14.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<3>.NEN
+ XI0.XI1.XI14.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<3>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<3>.MM_i_24 VDD! XI0.XI1.XI14.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<3>.MM_i_24_1 XI0.XI1.XI14.XI3<3>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<3>.MM_i_24_0 VDD! REG_DATA_2<3> XI0.XI1.XI14.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_2<3> XI0.XI1.XI14.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<3>.MM_i_24_1_48 XI0.XI1.XI14.XI3<3>.Y XI0.XI1.XI14.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<3>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<2>.MM_i_0 VSS! XI0.XI1.XI14.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<2>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<2>.MM_i_0_15 VSS! REG_DATA_2<2> XI0.XI1.XI14.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<2>.MM_i_0_15_63 XI0.XI1.XI14.XI3<2>.DUMMY1 REG_DATA_2<2>
+ XI0.XI1.XI14.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<2>.NEN
+ XI0.XI1.XI14.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<2>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<2>.MM_i_24 VDD! XI0.XI1.XI14.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<2>.MM_i_24_1 XI0.XI1.XI14.XI3<2>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<2>.MM_i_24_0 VDD! REG_DATA_2<2> XI0.XI1.XI14.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_2<2> XI0.XI1.XI14.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<2>.MM_i_24_1_48 XI0.XI1.XI14.XI3<2>.Y XI0.XI1.XI14.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<2>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<1>.MM_i_0 VSS! XI0.XI1.XI14.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<1>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<1>.MM_i_0_15 VSS! REG_DATA_2<1> XI0.XI1.XI14.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<1>.MM_i_0_15_63 XI0.XI1.XI14.XI3<1>.DUMMY1 REG_DATA_2<1>
+ XI0.XI1.XI14.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<1>.NEN
+ XI0.XI1.XI14.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<1>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<1>.MM_i_24 VDD! XI0.XI1.XI14.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<1>.MM_i_24_1 XI0.XI1.XI14.XI3<1>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<1>.MM_i_24_0 VDD! REG_DATA_2<1> XI0.XI1.XI14.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_2<1> XI0.XI1.XI14.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<1>.MM_i_24_1_48 XI0.XI1.XI14.XI3<1>.Y XI0.XI1.XI14.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<1>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<0>.MM_i_0 VSS! XI0.XI1.XI14.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<0>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<0>.MM_i_0_15 VSS! REG_DATA_2<0> XI0.XI1.XI14.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<0>.MM_i_0_15_63 XI0.XI1.XI14.XI3<0>.DUMMY1 REG_DATA_2<0>
+ XI0.XI1.XI14.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<0>.NEN
+ XI0.XI1.XI14.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<0>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<0>.MM_i_24 VDD! XI0.XI1.XI14.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<0>.MM_i_24_1 XI0.XI1.XI14.XI3<0>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<0>.MM_i_24_0 VDD! REG_DATA_2<0> XI0.XI1.XI14.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_2<0> XI0.XI1.XI14.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<0>.MM_i_24_1_48 XI0.XI1.XI14.XI3<0>.Y XI0.XI1.XI14.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<0>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<7>.MM_i_0 VSS! XI0.XI1.XI14.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<7>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<7>.MM_i_0_15 VSS! REG_DATA_2<7> XI0.XI1.XI14.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<7>.MM_i_0_15_63 XI0.XI1.XI14.XI3<7>.DUMMY1 REG_DATA_2<7>
+ XI0.XI1.XI14.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<7>.NEN
+ XI0.XI1.XI14.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<7>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<7>.MM_i_24 VDD! XI0.XI1.XI14.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<7>.MM_i_24_1 XI0.XI1.XI14.XI3<7>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<7>.MM_i_24_0 VDD! REG_DATA_2<7> XI0.XI1.XI14.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_2<7> XI0.XI1.XI14.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<7>.MM_i_24_1_48 XI0.XI1.XI14.XI3<7>.Y XI0.XI1.XI14.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<7>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<6>.MM_i_0 VSS! XI0.XI1.XI14.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<6>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<6>.MM_i_0_15 VSS! REG_DATA_2<6> XI0.XI1.XI14.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<6>.MM_i_0_15_63 XI0.XI1.XI14.XI3<6>.DUMMY1 REG_DATA_2<6>
+ XI0.XI1.XI14.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<6>.NEN
+ XI0.XI1.XI14.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<6>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<6>.MM_i_24 VDD! XI0.XI1.XI14.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<6>.MM_i_24_1 XI0.XI1.XI14.XI3<6>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<6>.MM_i_24_0 VDD! REG_DATA_2<6> XI0.XI1.XI14.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_2<6> XI0.XI1.XI14.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<6>.MM_i_24_1_48 XI0.XI1.XI14.XI3<6>.Y XI0.XI1.XI14.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<6>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<5>.MM_i_0 VSS! XI0.XI1.XI14.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<5>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<5>.MM_i_0_15 VSS! REG_DATA_2<5> XI0.XI1.XI14.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<5>.MM_i_0_15_63 XI0.XI1.XI14.XI3<5>.DUMMY1 REG_DATA_2<5>
+ XI0.XI1.XI14.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<5>.NEN
+ XI0.XI1.XI14.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<5>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<5>.MM_i_24 VDD! XI0.XI1.XI14.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<5>.MM_i_24_1 XI0.XI1.XI14.XI3<5>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<5>.MM_i_24_0 VDD! REG_DATA_2<5> XI0.XI1.XI14.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_2<5> XI0.XI1.XI14.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<5>.MM_i_24_1_48 XI0.XI1.XI14.XI3<5>.Y XI0.XI1.XI14.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<5>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<4>.MM_i_0 VSS! XI0.XI1.XI14.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<4>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<4>.MM_i_0_15 VSS! REG_DATA_2<4> XI0.XI1.XI14.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<4>.MM_i_0_15_63 XI0.XI1.XI14.XI3<4>.DUMMY1 REG_DATA_2<4>
+ XI0.XI1.XI14.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<4>.NEN
+ XI0.XI1.XI14.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<4>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<4>.MM_i_24 VDD! XI0.XI1.XI14.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<4>.MM_i_24_1 XI0.XI1.XI14.XI3<4>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<4>.MM_i_24_0 VDD! REG_DATA_2<4> XI0.XI1.XI14.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_2<4> XI0.XI1.XI14.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<4>.MM_i_24_1_48 XI0.XI1.XI14.XI3<4>.Y XI0.XI1.XI14.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<4>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<11>.MM_i_0 VSS! XI0.XI1.XI14.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<11>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<11>.MM_i_0_15 VSS! REG_DATA_2<11> XI0.XI1.XI14.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<11>.MM_i_0_15_63 XI0.XI1.XI14.XI3<11>.DUMMY1 REG_DATA_2<11>
+ XI0.XI1.XI14.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<11>.NEN
+ XI0.XI1.XI14.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<11>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<11>.MM_i_24 VDD! XI0.XI1.XI14.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<11>.MM_i_24_1 XI0.XI1.XI14.XI3<11>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<11>.MM_i_24_0 VDD! REG_DATA_2<11> XI0.XI1.XI14.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_2<11> XI0.XI1.XI14.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<11>.MM_i_24_1_48 XI0.XI1.XI14.XI3<11>.Y
+ XI0.XI1.XI14.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI14.XI3<11>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<10>.MM_i_0 VSS! XI0.XI1.XI14.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<10>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<10>.MM_i_0_15 VSS! REG_DATA_2<10> XI0.XI1.XI14.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<10>.MM_i_0_15_63 XI0.XI1.XI14.XI3<10>.DUMMY1 REG_DATA_2<10>
+ XI0.XI1.XI14.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<10>.NEN
+ XI0.XI1.XI14.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<10>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<10>.MM_i_24 VDD! XI0.XI1.XI14.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<10>.MM_i_24_1 XI0.XI1.XI14.XI3<10>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<10>.MM_i_24_0 VDD! REG_DATA_2<10> XI0.XI1.XI14.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_2<10> XI0.XI1.XI14.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<10>.MM_i_24_1_48 XI0.XI1.XI14.XI3<10>.Y
+ XI0.XI1.XI14.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI14.XI3<10>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<9>.MM_i_0 VSS! XI0.XI1.XI14.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<9>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<9>.MM_i_0_15 VSS! REG_DATA_2<9> XI0.XI1.XI14.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<9>.MM_i_0_15_63 XI0.XI1.XI14.XI3<9>.DUMMY1 REG_DATA_2<9>
+ XI0.XI1.XI14.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<9>.NEN
+ XI0.XI1.XI14.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<9>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<9>.MM_i_24 VDD! XI0.XI1.XI14.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<9>.MM_i_24_1 XI0.XI1.XI14.XI3<9>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<9>.MM_i_24_0 VDD! REG_DATA_2<9> XI0.XI1.XI14.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_2<9> XI0.XI1.XI14.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<9>.MM_i_24_1_48 XI0.XI1.XI14.XI3<9>.Y XI0.XI1.XI14.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<9>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<8>.MM_i_0 VSS! XI0.XI1.XI14.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<8>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<8>.MM_i_0_15 VSS! REG_DATA_2<8> XI0.XI1.XI14.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<8>.MM_i_0_15_63 XI0.XI1.XI14.XI3<8>.DUMMY1 REG_DATA_2<8>
+ XI0.XI1.XI14.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<8>.NEN
+ XI0.XI1.XI14.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<8>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<8>.MM_i_24 VDD! XI0.XI1.XI14.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<8>.MM_i_24_1 XI0.XI1.XI14.XI3<8>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<8>.MM_i_24_0 VDD! REG_DATA_2<8> XI0.XI1.XI14.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_2<8> XI0.XI1.XI14.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI14.XI3<8>.MM_i_24_1_48 XI0.XI1.XI14.XI3<8>.Y XI0.XI1.XI14.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI14.XI3<8>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<15>.MM_i_0 VSS! XI0.XI1.XI14.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<15>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<15>.MM_i_0_15 VSS! REG_DATA_2<15> XI0.XI1.XI14.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<15>.MM_i_0_15_63 XI0.XI1.XI14.XI3<15>.DUMMY1 REG_DATA_2<15>
+ XI0.XI1.XI14.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<15>.NEN
+ XI0.XI1.XI14.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<15>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<15>.MM_i_24 VDD! XI0.XI1.XI14.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<15>.MM_i_24_1 XI0.XI1.XI14.XI3<15>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<15>.MM_i_24_0 VDD! REG_DATA_2<15> XI0.XI1.XI14.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_2<15> XI0.XI1.XI14.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<15>.MM_i_24_1_48 XI0.XI1.XI14.XI3<15>.Y
+ XI0.XI1.XI14.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI14.XI3<15>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<14>.MM_i_0 VSS! XI0.XI1.XI14.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<14>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<14>.MM_i_0_15 VSS! REG_DATA_2<14> XI0.XI1.XI14.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<14>.MM_i_0_15_63 XI0.XI1.XI14.XI3<14>.DUMMY1 REG_DATA_2<14>
+ XI0.XI1.XI14.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<14>.NEN
+ XI0.XI1.XI14.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<14>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<14>.MM_i_24 VDD! XI0.XI1.XI14.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<14>.MM_i_24_1 XI0.XI1.XI14.XI3<14>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<14>.MM_i_24_0 VDD! REG_DATA_2<14> XI0.XI1.XI14.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_2<14> XI0.XI1.XI14.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<14>.MM_i_24_1_48 XI0.XI1.XI14.XI3<14>.Y
+ XI0.XI1.XI14.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI14.XI3<14>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<13>.MM_i_0 VSS! XI0.XI1.XI14.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<13>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<13>.MM_i_0_15 VSS! REG_DATA_2<13> XI0.XI1.XI14.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<13>.MM_i_0_15_63 XI0.XI1.XI14.XI3<13>.DUMMY1 REG_DATA_2<13>
+ XI0.XI1.XI14.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<13>.NEN
+ XI0.XI1.XI14.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<13>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<13>.MM_i_24 VDD! XI0.XI1.XI14.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<13>.MM_i_24_1 XI0.XI1.XI14.XI3<13>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<13>.MM_i_24_0 VDD! REG_DATA_2<13> XI0.XI1.XI14.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_2<13> XI0.XI1.XI14.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<13>.MM_i_24_1_48 XI0.XI1.XI14.XI3<13>.Y
+ XI0.XI1.XI14.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI14.XI3<13>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI14.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI14.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI14.XI3<12>.MM_i_0 VSS! XI0.XI1.XI14.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI14.XI3<12>.MM_i_0_14 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<12>.MM_i_0_15 VSS! REG_DATA_2<12> XI0.XI1.XI14.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<12>.MM_i_0_15_63 XI0.XI1.XI14.XI3<12>.DUMMY1 REG_DATA_2<12>
+ XI0.XI1.XI14.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI14.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI14.XI3<12>.NEN
+ XI0.XI1.XI14.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI14.XI3<12>.MM_i_17 VSS! XI0.NET1<10> XI0.XI1.XI14.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI14.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI14.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<12>.MM_i_24 VDD! XI0.XI1.XI14.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI14.XI3<12>.MM_i_24_1 XI0.XI1.XI14.XI3<12>.DUMMY0 XI0.NET1<10>
+ XI0.XI1.XI14.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI14.XI3<12>.MM_i_24_0 VDD! REG_DATA_2<12> XI0.XI1.XI14.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_2<12> XI0.XI1.XI14.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI14.XI3<12>.MM_i_24_1_48 XI0.XI1.XI14.XI3<12>.Y
+ XI0.XI1.XI14.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI14.XI3<12>.MM_i_42 VDD! XI0.NET1<10> XI0.XI1.XI14.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<3>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<3>.MM_i_0 VSS! XI0.XI1.XI13.XI3<3>.X RD_DATA_0<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<3>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<3>.MM_i_0_15 VSS! REG_DATA_1<3> XI0.XI1.XI13.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<3>.MM_i_0_15_63 XI0.XI1.XI13.XI3<3>.DUMMY1 REG_DATA_1<3>
+ XI0.XI1.XI13.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<3>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<3>.NEN
+ XI0.XI1.XI13.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<3>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<3>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<3>.MM_i_24 VDD! XI0.XI1.XI13.XI3<3>.Y RD_DATA_0<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<3>.MM_i_24_1 XI0.XI1.XI13.XI3<3>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<3>.MM_i_24_0 VDD! REG_DATA_1<3> XI0.XI1.XI13.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_1<3> XI0.XI1.XI13.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<3>.MM_i_24_1_48 XI0.XI1.XI13.XI3<3>.Y XI0.XI1.XI13.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<3>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<2>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<2>.MM_i_0 VSS! XI0.XI1.XI13.XI3<2>.X RD_DATA_0<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<2>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<2>.MM_i_0_15 VSS! REG_DATA_1<2> XI0.XI1.XI13.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<2>.MM_i_0_15_63 XI0.XI1.XI13.XI3<2>.DUMMY1 REG_DATA_1<2>
+ XI0.XI1.XI13.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<2>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<2>.NEN
+ XI0.XI1.XI13.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<2>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<2>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<2>.MM_i_24 VDD! XI0.XI1.XI13.XI3<2>.Y RD_DATA_0<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<2>.MM_i_24_1 XI0.XI1.XI13.XI3<2>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<2>.MM_i_24_0 VDD! REG_DATA_1<2> XI0.XI1.XI13.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_1<2> XI0.XI1.XI13.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<2>.MM_i_24_1_48 XI0.XI1.XI13.XI3<2>.Y XI0.XI1.XI13.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<2>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<1>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<1>.MM_i_0 VSS! XI0.XI1.XI13.XI3<1>.X RD_DATA_0<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<1>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<1>.MM_i_0_15 VSS! REG_DATA_1<1> XI0.XI1.XI13.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<1>.MM_i_0_15_63 XI0.XI1.XI13.XI3<1>.DUMMY1 REG_DATA_1<1>
+ XI0.XI1.XI13.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<1>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<1>.NEN
+ XI0.XI1.XI13.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<1>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<1>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<1>.MM_i_24 VDD! XI0.XI1.XI13.XI3<1>.Y RD_DATA_0<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<1>.MM_i_24_1 XI0.XI1.XI13.XI3<1>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<1>.MM_i_24_0 VDD! REG_DATA_1<1> XI0.XI1.XI13.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_1<1> XI0.XI1.XI13.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<1>.MM_i_24_1_48 XI0.XI1.XI13.XI3<1>.Y XI0.XI1.XI13.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<1>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<0>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<0>.MM_i_0 VSS! XI0.XI1.XI13.XI3<0>.X RD_DATA_0<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<0>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<0>.MM_i_0_15 VSS! REG_DATA_1<0> XI0.XI1.XI13.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<0>.MM_i_0_15_63 XI0.XI1.XI13.XI3<0>.DUMMY1 REG_DATA_1<0>
+ XI0.XI1.XI13.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<0>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<0>.NEN
+ XI0.XI1.XI13.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<0>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<0>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<0>.MM_i_24 VDD! XI0.XI1.XI13.XI3<0>.Y RD_DATA_0<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<0>.MM_i_24_1 XI0.XI1.XI13.XI3<0>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<0>.MM_i_24_0 VDD! REG_DATA_1<0> XI0.XI1.XI13.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_1<0> XI0.XI1.XI13.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<0>.MM_i_24_1_48 XI0.XI1.XI13.XI3<0>.Y XI0.XI1.XI13.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<0>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<7>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<7>.MM_i_0 VSS! XI0.XI1.XI13.XI3<7>.X RD_DATA_0<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<7>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<7>.MM_i_0_15 VSS! REG_DATA_1<7> XI0.XI1.XI13.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<7>.MM_i_0_15_63 XI0.XI1.XI13.XI3<7>.DUMMY1 REG_DATA_1<7>
+ XI0.XI1.XI13.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<7>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<7>.NEN
+ XI0.XI1.XI13.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<7>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<7>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<7>.MM_i_24 VDD! XI0.XI1.XI13.XI3<7>.Y RD_DATA_0<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<7>.MM_i_24_1 XI0.XI1.XI13.XI3<7>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<7>.MM_i_24_0 VDD! REG_DATA_1<7> XI0.XI1.XI13.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_1<7> XI0.XI1.XI13.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<7>.MM_i_24_1_48 XI0.XI1.XI13.XI3<7>.Y XI0.XI1.XI13.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<7>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<6>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<6>.MM_i_0 VSS! XI0.XI1.XI13.XI3<6>.X RD_DATA_0<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<6>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<6>.MM_i_0_15 VSS! REG_DATA_1<6> XI0.XI1.XI13.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<6>.MM_i_0_15_63 XI0.XI1.XI13.XI3<6>.DUMMY1 REG_DATA_1<6>
+ XI0.XI1.XI13.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<6>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<6>.NEN
+ XI0.XI1.XI13.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<6>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<6>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<6>.MM_i_24 VDD! XI0.XI1.XI13.XI3<6>.Y RD_DATA_0<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<6>.MM_i_24_1 XI0.XI1.XI13.XI3<6>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<6>.MM_i_24_0 VDD! REG_DATA_1<6> XI0.XI1.XI13.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_1<6> XI0.XI1.XI13.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<6>.MM_i_24_1_48 XI0.XI1.XI13.XI3<6>.Y XI0.XI1.XI13.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<6>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<5>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<5>.MM_i_0 VSS! XI0.XI1.XI13.XI3<5>.X RD_DATA_0<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<5>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<5>.MM_i_0_15 VSS! REG_DATA_1<5> XI0.XI1.XI13.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<5>.MM_i_0_15_63 XI0.XI1.XI13.XI3<5>.DUMMY1 REG_DATA_1<5>
+ XI0.XI1.XI13.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<5>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<5>.NEN
+ XI0.XI1.XI13.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<5>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<5>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<5>.MM_i_24 VDD! XI0.XI1.XI13.XI3<5>.Y RD_DATA_0<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<5>.MM_i_24_1 XI0.XI1.XI13.XI3<5>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<5>.MM_i_24_0 VDD! REG_DATA_1<5> XI0.XI1.XI13.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_1<5> XI0.XI1.XI13.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<5>.MM_i_24_1_48 XI0.XI1.XI13.XI3<5>.Y XI0.XI1.XI13.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<5>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<4>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<4>.MM_i_0 VSS! XI0.XI1.XI13.XI3<4>.X RD_DATA_0<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<4>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<4>.MM_i_0_15 VSS! REG_DATA_1<4> XI0.XI1.XI13.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<4>.MM_i_0_15_63 XI0.XI1.XI13.XI3<4>.DUMMY1 REG_DATA_1<4>
+ XI0.XI1.XI13.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<4>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<4>.NEN
+ XI0.XI1.XI13.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<4>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<4>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<4>.MM_i_24 VDD! XI0.XI1.XI13.XI3<4>.Y RD_DATA_0<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<4>.MM_i_24_1 XI0.XI1.XI13.XI3<4>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<4>.MM_i_24_0 VDD! REG_DATA_1<4> XI0.XI1.XI13.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_1<4> XI0.XI1.XI13.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<4>.MM_i_24_1_48 XI0.XI1.XI13.XI3<4>.Y XI0.XI1.XI13.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<4>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<11>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<11>.MM_i_0 VSS! XI0.XI1.XI13.XI3<11>.X RD_DATA_0<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<11>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<11>.MM_i_0_15 VSS! REG_DATA_1<11> XI0.XI1.XI13.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<11>.MM_i_0_15_63 XI0.XI1.XI13.XI3<11>.DUMMY1 REG_DATA_1<11>
+ XI0.XI1.XI13.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<11>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<11>.NEN
+ XI0.XI1.XI13.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<11>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<11>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<11>.MM_i_24 VDD! XI0.XI1.XI13.XI3<11>.Y RD_DATA_0<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<11>.MM_i_24_1 XI0.XI1.XI13.XI3<11>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<11>.MM_i_24_0 VDD! REG_DATA_1<11> XI0.XI1.XI13.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_1<11> XI0.XI1.XI13.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<11>.MM_i_24_1_48 XI0.XI1.XI13.XI3<11>.Y
+ XI0.XI1.XI13.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI13.XI3<11>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<10>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<10>.MM_i_0 VSS! XI0.XI1.XI13.XI3<10>.X RD_DATA_0<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<10>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<10>.MM_i_0_15 VSS! REG_DATA_1<10> XI0.XI1.XI13.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<10>.MM_i_0_15_63 XI0.XI1.XI13.XI3<10>.DUMMY1 REG_DATA_1<10>
+ XI0.XI1.XI13.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<10>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<10>.NEN
+ XI0.XI1.XI13.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<10>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<10>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<10>.MM_i_24 VDD! XI0.XI1.XI13.XI3<10>.Y RD_DATA_0<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<10>.MM_i_24_1 XI0.XI1.XI13.XI3<10>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<10>.MM_i_24_0 VDD! REG_DATA_1<10> XI0.XI1.XI13.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_1<10> XI0.XI1.XI13.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<10>.MM_i_24_1_48 XI0.XI1.XI13.XI3<10>.Y
+ XI0.XI1.XI13.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI13.XI3<10>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<9>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<9>.MM_i_0 VSS! XI0.XI1.XI13.XI3<9>.X RD_DATA_0<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<9>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<9>.MM_i_0_15 VSS! REG_DATA_1<9> XI0.XI1.XI13.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<9>.MM_i_0_15_63 XI0.XI1.XI13.XI3<9>.DUMMY1 REG_DATA_1<9>
+ XI0.XI1.XI13.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<9>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<9>.NEN
+ XI0.XI1.XI13.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<9>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<9>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<9>.MM_i_24 VDD! XI0.XI1.XI13.XI3<9>.Y RD_DATA_0<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<9>.MM_i_24_1 XI0.XI1.XI13.XI3<9>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<9>.MM_i_24_0 VDD! REG_DATA_1<9> XI0.XI1.XI13.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_1<9> XI0.XI1.XI13.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<9>.MM_i_24_1_48 XI0.XI1.XI13.XI3<9>.Y XI0.XI1.XI13.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<9>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<8>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<8>.MM_i_0 VSS! XI0.XI1.XI13.XI3<8>.X RD_DATA_0<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<8>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<8>.MM_i_0_15 VSS! REG_DATA_1<8> XI0.XI1.XI13.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<8>.MM_i_0_15_63 XI0.XI1.XI13.XI3<8>.DUMMY1 REG_DATA_1<8>
+ XI0.XI1.XI13.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<8>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<8>.NEN
+ XI0.XI1.XI13.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<8>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<8>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<8>.MM_i_24 VDD! XI0.XI1.XI13.XI3<8>.Y RD_DATA_0<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<8>.MM_i_24_1 XI0.XI1.XI13.XI3<8>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<8>.MM_i_24_0 VDD! REG_DATA_1<8> XI0.XI1.XI13.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_1<8> XI0.XI1.XI13.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI0.XI1.XI13.XI3<8>.MM_i_24_1_48 XI0.XI1.XI13.XI3<8>.Y XI0.XI1.XI13.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI0.XI1.XI13.XI3<8>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<15>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<15>.MM_i_0 VSS! XI0.XI1.XI13.XI3<15>.X RD_DATA_0<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<15>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<15>.MM_i_0_15 VSS! REG_DATA_1<15> XI0.XI1.XI13.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<15>.MM_i_0_15_63 XI0.XI1.XI13.XI3<15>.DUMMY1 REG_DATA_1<15>
+ XI0.XI1.XI13.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<15>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<15>.NEN
+ XI0.XI1.XI13.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<15>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<15>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<15>.MM_i_24 VDD! XI0.XI1.XI13.XI3<15>.Y RD_DATA_0<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<15>.MM_i_24_1 XI0.XI1.XI13.XI3<15>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<15>.MM_i_24_0 VDD! REG_DATA_1<15> XI0.XI1.XI13.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_1<15> XI0.XI1.XI13.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<15>.MM_i_24_1_48 XI0.XI1.XI13.XI3<15>.Y
+ XI0.XI1.XI13.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI13.XI3<15>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<14>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<14>.MM_i_0 VSS! XI0.XI1.XI13.XI3<14>.X RD_DATA_0<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<14>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<14>.MM_i_0_15 VSS! REG_DATA_1<14> XI0.XI1.XI13.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<14>.MM_i_0_15_63 XI0.XI1.XI13.XI3<14>.DUMMY1 REG_DATA_1<14>
+ XI0.XI1.XI13.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<14>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<14>.NEN
+ XI0.XI1.XI13.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<14>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<14>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<14>.MM_i_24 VDD! XI0.XI1.XI13.XI3<14>.Y RD_DATA_0<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<14>.MM_i_24_1 XI0.XI1.XI13.XI3<14>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<14>.MM_i_24_0 VDD! REG_DATA_1<14> XI0.XI1.XI13.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_1<14> XI0.XI1.XI13.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<14>.MM_i_24_1_48 XI0.XI1.XI13.XI3<14>.Y
+ XI0.XI1.XI13.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI13.XI3<14>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<13>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<13>.MM_i_0 VSS! XI0.XI1.XI13.XI3<13>.X RD_DATA_0<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<13>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<13>.MM_i_0_15 VSS! REG_DATA_1<13> XI0.XI1.XI13.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<13>.MM_i_0_15_63 XI0.XI1.XI13.XI3<13>.DUMMY1 REG_DATA_1<13>
+ XI0.XI1.XI13.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<13>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<13>.NEN
+ XI0.XI1.XI13.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<13>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<13>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<13>.MM_i_24 VDD! XI0.XI1.XI13.XI3<13>.Y RD_DATA_0<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<13>.MM_i_24_1 XI0.XI1.XI13.XI3<13>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<13>.MM_i_24_0 VDD! REG_DATA_1<13> XI0.XI1.XI13.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_1<13> XI0.XI1.XI13.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<13>.MM_i_24_1_48 XI0.XI1.XI13.XI3<13>.Y
+ XI0.XI1.XI13.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI13.XI3<13>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI0.XI1.XI13.XI3<12>.MM_i_0_6 VSS! XI0.XI1.XI13.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI0.XI1.XI13.XI3<12>.MM_i_0 VSS! XI0.XI1.XI13.XI3<12>.X RD_DATA_0<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI0.XI1.XI13.XI3<12>.MM_i_0_14 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<12>.MM_i_0_15 VSS! REG_DATA_1<12> XI0.XI1.XI13.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<12>.MM_i_0_15_63 XI0.XI1.XI13.XI3<12>.DUMMY1 REG_DATA_1<12>
+ XI0.XI1.XI13.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI0.XI1.XI13.XI3<12>.MM_i_0_14_47 VSS! XI0.XI1.XI13.XI3<12>.NEN
+ XI0.XI1.XI13.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI0.XI1.XI13.XI3<12>.MM_i_17 VSS! XI0.NET1<11> XI0.XI1.XI13.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI0.XI1.XI13.XI3<12>.MM_i_24_3 VDD! XI0.XI1.XI13.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<12>.MM_i_24 VDD! XI0.XI1.XI13.XI3<12>.Y RD_DATA_0<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI0.XI1.XI13.XI3<12>.MM_i_24_1 XI0.XI1.XI13.XI3<12>.DUMMY0 XI0.NET1<11>
+ XI0.XI1.XI13.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI0.XI1.XI13.XI3<12>.MM_i_24_0 VDD! REG_DATA_1<12> XI0.XI1.XI13.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_1<12> XI0.XI1.XI13.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI0.XI1.XI13.XI3<12>.MM_i_24_1_48 XI0.XI1.XI13.XI3<12>.Y
+ XI0.XI1.XI13.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI0.XI1.XI13.XI3<12>.MM_i_42 VDD! XI0.NET1<11> XI0.XI1.XI13.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI0.XI24.MM_i_1 XI2.XI0.XI24.NET_0 XI2.XI0.NET_11XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI24.MM_i_0 XI2.NET1<0> XI2.XI0.NET_XX00 XI2.XI0.XI24.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI24.MM_i_3 XI2.NET1<0> XI2.XI0.NET_11XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI24.MM_i_2 VDD! XI2.XI0.NET_XX00 XI2.NET1<0> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI23.MM_i_1 XI2.XI0.XI23.NET_0 XI2.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI23.MM_i_0 XI2.NET1<1> XI2.XI0.NET_XX11 XI2.XI0.XI23.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI23.MM_i_3 XI2.NET1<1> XI2.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI23.MM_i_2 VDD! XI2.XI0.NET_XX11 XI2.NET1<1> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI22.MM_i_1 XI2.XI0.XI22.NET_0 XI2.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI22.MM_i_0 XI2.NET1<2> XI2.XI0.NET_XX10 XI2.XI0.XI22.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI22.MM_i_3 XI2.NET1<2> XI2.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI22.MM_i_2 VDD! XI2.XI0.NET_XX10 XI2.NET1<2> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI21.MM_i_1 XI2.XI0.XI21.NET_0 XI2.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI21.MM_i_0 XI2.NET1<3> XI2.XI0.NET_XX01 XI2.XI0.XI21.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI21.MM_i_3 XI2.NET1<3> XI2.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI21.MM_i_2 VDD! XI2.XI0.NET_XX01 XI2.NET1<3> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI20.MM_i_1 XI2.XI0.XI20.NET_0 XI2.XI0.NET_10XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI20.MM_i_0 XI2.NET1<4> XI2.XI0.NET_XX00 XI2.XI0.XI20.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI20.MM_i_3 XI2.NET1<4> XI2.XI0.NET_10XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI20.MM_i_2 VDD! XI2.XI0.NET_XX00 XI2.NET1<4> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI19.MM_i_1 XI2.XI0.XI19.NET_0 XI2.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI19.MM_i_0 XI2.NET1<5> XI2.XI0.NET_XX11 XI2.XI0.XI19.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI19.MM_i_3 XI2.NET1<5> XI2.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI19.MM_i_2 VDD! XI2.XI0.NET_XX11 XI2.NET1<5> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI18.MM_i_1 XI2.XI0.XI18.NET_0 XI2.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI18.MM_i_0 XI2.NET1<6> XI2.XI0.NET_XX10 XI2.XI0.XI18.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI18.MM_i_3 XI2.NET1<6> XI2.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI18.MM_i_2 VDD! XI2.XI0.NET_XX10 XI2.NET1<6> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI17.MM_i_1 XI2.XI0.XI17.NET_0 XI2.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI17.MM_i_0 XI2.NET1<7> XI2.XI0.NET_XX01 XI2.XI0.XI17.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI17.MM_i_3 XI2.NET1<7> XI2.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI17.MM_i_2 VDD! XI2.XI0.NET_XX01 XI2.NET1<7> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI16.MM_i_1 XI2.XI0.XI16.NET_0 XI2.XI0.NET_01XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI16.MM_i_0 XI2.NET1<8> XI2.XI0.NET_XX00 XI2.XI0.XI16.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI16.MM_i_3 XI2.NET1<8> XI2.XI0.NET_01XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI16.MM_i_2 VDD! XI2.XI0.NET_XX00 XI2.NET1<8> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI15.MM_i_1 XI2.XI0.XI15.NET_0 XI2.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI15.MM_i_0 XI2.NET1<9> XI2.XI0.NET_XX11 XI2.XI0.XI15.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI15.MM_i_3 XI2.NET1<9> XI2.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI15.MM_i_2 VDD! XI2.XI0.NET_XX11 XI2.NET1<9> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI14.MM_i_1 XI2.XI0.XI14.NET_0 XI2.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI14.MM_i_0 XI2.NET1<10> XI2.XI0.NET_XX10 XI2.XI0.XI14.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI14.MM_i_3 XI2.NET1<10> XI2.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI14.MM_i_2 VDD! XI2.XI0.NET_XX10 XI2.NET1<10> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI13.MM_i_1 XI2.XI0.XI13.NET_0 XI2.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI13.MM_i_0 XI2.NET1<11> XI2.XI0.NET_XX01 XI2.XI0.XI13.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI13.MM_i_3 XI2.NET1<11> XI2.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI13.MM_i_2 VDD! XI2.XI0.NET_XX01 XI2.NET1<11> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI12.MM_i_1 XI2.XI0.XI12.NET_0 XI2.XI0.NET_00XX VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI0.XI12.MM_i_0 XI2.NET1<12> XI2.XI0.NET_XX00 XI2.XI0.XI12.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI12.MM_i_3 XI2.NET1<12> XI2.XI0.NET_00XX VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI0.XI12.MM_i_2 VDD! XI2.XI0.NET_XX00 XI2.NET1<12> VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI11.MM_i_2 XI2.XI0.XI11.NET_0 RD_ADDR_1<2> XI2.XI0.XI11.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI11.MM_i_3 VSS! RD_ADDR_1<3> XI2.XI0.XI11.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI11.MM_i_0 XI2.XI0.NET_11XX XI2.XI0.XI11.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI11.MM_i_4 XI2.XI0.XI11.ZN_NEG RD_ADDR_1<2> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI11.MM_i_5 VDD! RD_ADDR_1<3> XI2.XI0.XI11.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI11.MM_i_1 XI2.XI0.NET_11XX XI2.XI0.XI11.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI7.MM_i_2 XI2.XI0.XI7.NET_0 RD_ADDR_1<0> XI2.XI0.XI7.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI7.MM_i_3 VSS! RD_ADDR_1<1> XI2.XI0.XI7.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI7.MM_i_0 XI2.XI0.NET_XX11 XI2.XI0.XI7.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI7.MM_i_4 XI2.XI0.XI7.ZN_NEG RD_ADDR_1<0> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI7.MM_i_5 VDD! RD_ADDR_1<1> XI2.XI0.XI7.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI7.MM_i_1 XI2.XI0.NET_XX11 XI2.XI0.XI7.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI10.MM_i_2 XI2.XI0.XI10.NET_0 XI2.XI0.ADDR_BAR<2> XI2.XI0.XI10.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI10.MM_i_3 VSS! RD_ADDR_1<3> XI2.XI0.XI10.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI10.MM_i_0 XI2.XI0.NET_10XX XI2.XI0.XI10.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI10.MM_i_4 XI2.XI0.XI10.ZN_NEG XI2.XI0.ADDR_BAR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI10.MM_i_5 VDD! RD_ADDR_1<3> XI2.XI0.XI10.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI10.MM_i_1 XI2.XI0.NET_10XX XI2.XI0.XI10.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI6.MM_i_2 XI2.XI0.XI6.NET_0 XI2.XI0.ADDR_BAR<0> XI2.XI0.XI6.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI6.MM_i_3 VSS! RD_ADDR_1<1> XI2.XI0.XI6.NET_0 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI6.MM_i_0 XI2.XI0.NET_XX10 XI2.XI0.XI6.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI6.MM_i_4 XI2.XI0.XI6.ZN_NEG XI2.XI0.ADDR_BAR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI6.MM_i_5 VDD! RD_ADDR_1<1> XI2.XI0.XI6.ZN_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI6.MM_i_1 XI2.XI0.NET_XX10 XI2.XI0.XI6.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI9.MM_i_2 XI2.XI0.XI9.NET_0 RD_ADDR_1<2> XI2.XI0.XI9.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI9.MM_i_3 VSS! XI2.XI0.ADDR_BAR<3> XI2.XI0.XI9.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI9.MM_i_0 XI2.XI0.NET_01XX XI2.XI0.XI9.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI9.MM_i_4 XI2.XI0.XI9.ZN_NEG RD_ADDR_1<2> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI9.MM_i_5 VDD! XI2.XI0.ADDR_BAR<3> XI2.XI0.XI9.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI9.MM_i_1 XI2.XI0.NET_01XX XI2.XI0.XI9.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI5.MM_i_2 XI2.XI0.XI5.NET_0 RD_ADDR_1<0> XI2.XI0.XI5.ZN_NEG VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI5.MM_i_3 VSS! XI2.XI0.ADDR_BAR<1> XI2.XI0.XI5.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI5.MM_i_0 XI2.XI0.NET_XX01 XI2.XI0.XI5.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI5.MM_i_4 XI2.XI0.XI5.ZN_NEG RD_ADDR_1<0> VDD! VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI5.MM_i_5 VDD! XI2.XI0.ADDR_BAR<1> XI2.XI0.XI5.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI5.MM_i_1 XI2.XI0.NET_XX01 XI2.XI0.XI5.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI8.MM_i_2 XI2.XI0.XI8.NET_0 XI2.XI0.ADDR_BAR<2> XI2.XI0.XI8.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI8.MM_i_3 VSS! XI2.XI0.ADDR_BAR<3> XI2.XI0.XI8.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI8.MM_i_0 XI2.XI0.NET_00XX XI2.XI0.XI8.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI8.MM_i_4 XI2.XI0.XI8.ZN_NEG XI2.XI0.ADDR_BAR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI8.MM_i_5 VDD! XI2.XI0.ADDR_BAR<3> XI2.XI0.XI8.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI8.MM_i_1 XI2.XI0.NET_00XX XI2.XI0.XI8.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI4.MM_i_2 XI2.XI0.XI4.NET_0 XI2.XI0.ADDR_BAR<0> XI2.XI0.XI4.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI2.XI0.XI4.MM_i_3 VSS! XI2.XI0.ADDR_BAR<1> XI2.XI0.XI4.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI2.XI0.XI4.MM_i_0 XI2.XI0.NET_XX00 XI2.XI0.XI4.ZN_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI0.XI4.MM_i_4 XI2.XI0.XI4.ZN_NEG XI2.XI0.ADDR_BAR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI2.XI0.XI4.MM_i_5 VDD! XI2.XI0.ADDR_BAR<1> XI2.XI0.XI4.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI2.XI0.XI4.MM_i_1 XI2.XI0.NET_XX00 XI2.XI0.XI4.ZN_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI2.XI0.XI2.MM_i_0 XI2.XI0.ADDR_BAR<2> RD_ADDR_1<2> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI2.XI0.XI2.MM_i_1 XI2.XI0.ADDR_BAR<2> RD_ADDR_1<2> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI2.XI0.XI0.MM_i_0 XI2.XI0.ADDR_BAR<0> RD_ADDR_1<0> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI2.XI0.XI0.MM_i_1 XI2.XI0.ADDR_BAR<0> RD_ADDR_1<0> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI2.XI0.XI3.MM_i_0 XI2.XI0.ADDR_BAR<3> RD_ADDR_1<3> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI2.XI0.XI3.MM_i_1 XI2.XI0.ADDR_BAR<3> RD_ADDR_1<3> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI2.XI0.XI1.MM_i_0 XI2.XI0.ADDR_BAR<1> RD_ADDR_1<1> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI2.XI0.XI1.MM_i_1 XI2.XI0.ADDR_BAR<1> RD_ADDR_1<1> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<3>.MM_i_0 VSS! XI2.XI1.XI15.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<3>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<3>.MM_i_0_15 VSS! REG_DATA_0<3> XI2.XI1.XI15.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<3>.MM_i_0_15_63 XI2.XI1.XI15.XI3<3>.DUMMY1 REG_DATA_0<3>
+ XI2.XI1.XI15.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<3>.NEN
+ XI2.XI1.XI15.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<3>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<3>.MM_i_24 VDD! XI2.XI1.XI15.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<3>.MM_i_24_1 XI2.XI1.XI15.XI3<3>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<3>.MM_i_24_0 VDD! REG_DATA_0<3> XI2.XI1.XI15.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_0<3> XI2.XI1.XI15.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<3>.MM_i_24_1_48 XI2.XI1.XI15.XI3<3>.Y XI2.XI1.XI15.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<3>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<2>.MM_i_0 VSS! XI2.XI1.XI15.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<2>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<2>.MM_i_0_15 VSS! REG_DATA_0<2> XI2.XI1.XI15.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<2>.MM_i_0_15_63 XI2.XI1.XI15.XI3<2>.DUMMY1 REG_DATA_0<2>
+ XI2.XI1.XI15.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<2>.NEN
+ XI2.XI1.XI15.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<2>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<2>.MM_i_24 VDD! XI2.XI1.XI15.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<2>.MM_i_24_1 XI2.XI1.XI15.XI3<2>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<2>.MM_i_24_0 VDD! REG_DATA_0<2> XI2.XI1.XI15.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_0<2> XI2.XI1.XI15.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<2>.MM_i_24_1_48 XI2.XI1.XI15.XI3<2>.Y XI2.XI1.XI15.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<2>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<1>.MM_i_0 VSS! XI2.XI1.XI15.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<1>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<1>.MM_i_0_15 VSS! REG_DATA_0<1> XI2.XI1.XI15.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<1>.MM_i_0_15_63 XI2.XI1.XI15.XI3<1>.DUMMY1 REG_DATA_0<1>
+ XI2.XI1.XI15.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<1>.NEN
+ XI2.XI1.XI15.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<1>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<1>.MM_i_24 VDD! XI2.XI1.XI15.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<1>.MM_i_24_1 XI2.XI1.XI15.XI3<1>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<1>.MM_i_24_0 VDD! REG_DATA_0<1> XI2.XI1.XI15.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_0<1> XI2.XI1.XI15.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<1>.MM_i_24_1_48 XI2.XI1.XI15.XI3<1>.Y XI2.XI1.XI15.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<1>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<0>.MM_i_0 VSS! XI2.XI1.XI15.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<0>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<0>.MM_i_0_15 VSS! REG_DATA_0<0> XI2.XI1.XI15.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<0>.MM_i_0_15_63 XI2.XI1.XI15.XI3<0>.DUMMY1 REG_DATA_0<0>
+ XI2.XI1.XI15.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<0>.NEN
+ XI2.XI1.XI15.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<0>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<0>.MM_i_24 VDD! XI2.XI1.XI15.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<0>.MM_i_24_1 XI2.XI1.XI15.XI3<0>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<0>.MM_i_24_0 VDD! REG_DATA_0<0> XI2.XI1.XI15.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_0<0> XI2.XI1.XI15.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<0>.MM_i_24_1_48 XI2.XI1.XI15.XI3<0>.Y XI2.XI1.XI15.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<0>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<7>.MM_i_0 VSS! XI2.XI1.XI15.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<7>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<7>.MM_i_0_15 VSS! REG_DATA_0<7> XI2.XI1.XI15.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<7>.MM_i_0_15_63 XI2.XI1.XI15.XI3<7>.DUMMY1 REG_DATA_0<7>
+ XI2.XI1.XI15.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<7>.NEN
+ XI2.XI1.XI15.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<7>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<7>.MM_i_24 VDD! XI2.XI1.XI15.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<7>.MM_i_24_1 XI2.XI1.XI15.XI3<7>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<7>.MM_i_24_0 VDD! REG_DATA_0<7> XI2.XI1.XI15.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_0<7> XI2.XI1.XI15.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<7>.MM_i_24_1_48 XI2.XI1.XI15.XI3<7>.Y XI2.XI1.XI15.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<7>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<6>.MM_i_0 VSS! XI2.XI1.XI15.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<6>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<6>.MM_i_0_15 VSS! REG_DATA_0<6> XI2.XI1.XI15.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<6>.MM_i_0_15_63 XI2.XI1.XI15.XI3<6>.DUMMY1 REG_DATA_0<6>
+ XI2.XI1.XI15.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<6>.NEN
+ XI2.XI1.XI15.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<6>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<6>.MM_i_24 VDD! XI2.XI1.XI15.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<6>.MM_i_24_1 XI2.XI1.XI15.XI3<6>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<6>.MM_i_24_0 VDD! REG_DATA_0<6> XI2.XI1.XI15.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_0<6> XI2.XI1.XI15.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<6>.MM_i_24_1_48 XI2.XI1.XI15.XI3<6>.Y XI2.XI1.XI15.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<6>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<5>.MM_i_0 VSS! XI2.XI1.XI15.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<5>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<5>.MM_i_0_15 VSS! REG_DATA_0<5> XI2.XI1.XI15.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<5>.MM_i_0_15_63 XI2.XI1.XI15.XI3<5>.DUMMY1 REG_DATA_0<5>
+ XI2.XI1.XI15.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<5>.NEN
+ XI2.XI1.XI15.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<5>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<5>.MM_i_24 VDD! XI2.XI1.XI15.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<5>.MM_i_24_1 XI2.XI1.XI15.XI3<5>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<5>.MM_i_24_0 VDD! REG_DATA_0<5> XI2.XI1.XI15.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_0<5> XI2.XI1.XI15.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<5>.MM_i_24_1_48 XI2.XI1.XI15.XI3<5>.Y XI2.XI1.XI15.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<5>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<4>.MM_i_0 VSS! XI2.XI1.XI15.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<4>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<4>.MM_i_0_15 VSS! REG_DATA_0<4> XI2.XI1.XI15.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<4>.MM_i_0_15_63 XI2.XI1.XI15.XI3<4>.DUMMY1 REG_DATA_0<4>
+ XI2.XI1.XI15.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<4>.NEN
+ XI2.XI1.XI15.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<4>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<4>.MM_i_24 VDD! XI2.XI1.XI15.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<4>.MM_i_24_1 XI2.XI1.XI15.XI3<4>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<4>.MM_i_24_0 VDD! REG_DATA_0<4> XI2.XI1.XI15.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_0<4> XI2.XI1.XI15.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<4>.MM_i_24_1_48 XI2.XI1.XI15.XI3<4>.Y XI2.XI1.XI15.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<4>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<11>.MM_i_0 VSS! XI2.XI1.XI15.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<11>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<11>.MM_i_0_15 VSS! REG_DATA_0<11> XI2.XI1.XI15.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<11>.MM_i_0_15_63 XI2.XI1.XI15.XI3<11>.DUMMY1 REG_DATA_0<11>
+ XI2.XI1.XI15.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<11>.NEN
+ XI2.XI1.XI15.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<11>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<11>.MM_i_24 VDD! XI2.XI1.XI15.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<11>.MM_i_24_1 XI2.XI1.XI15.XI3<11>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<11>.MM_i_24_0 VDD! REG_DATA_0<11> XI2.XI1.XI15.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_0<11> XI2.XI1.XI15.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<11>.MM_i_24_1_48 XI2.XI1.XI15.XI3<11>.Y
+ XI2.XI1.XI15.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI15.XI3<11>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<10>.MM_i_0 VSS! XI2.XI1.XI15.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<10>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<10>.MM_i_0_15 VSS! REG_DATA_0<10> XI2.XI1.XI15.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<10>.MM_i_0_15_63 XI2.XI1.XI15.XI3<10>.DUMMY1 REG_DATA_0<10>
+ XI2.XI1.XI15.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<10>.NEN
+ XI2.XI1.XI15.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<10>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<10>.MM_i_24 VDD! XI2.XI1.XI15.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<10>.MM_i_24_1 XI2.XI1.XI15.XI3<10>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<10>.MM_i_24_0 VDD! REG_DATA_0<10> XI2.XI1.XI15.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_0<10> XI2.XI1.XI15.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<10>.MM_i_24_1_48 XI2.XI1.XI15.XI3<10>.Y
+ XI2.XI1.XI15.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI15.XI3<10>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<9>.MM_i_0 VSS! XI2.XI1.XI15.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<9>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<9>.MM_i_0_15 VSS! REG_DATA_0<9> XI2.XI1.XI15.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<9>.MM_i_0_15_63 XI2.XI1.XI15.XI3<9>.DUMMY1 REG_DATA_0<9>
+ XI2.XI1.XI15.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<9>.NEN
+ XI2.XI1.XI15.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<9>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<9>.MM_i_24 VDD! XI2.XI1.XI15.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<9>.MM_i_24_1 XI2.XI1.XI15.XI3<9>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<9>.MM_i_24_0 VDD! REG_DATA_0<9> XI2.XI1.XI15.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_0<9> XI2.XI1.XI15.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<9>.MM_i_24_1_48 XI2.XI1.XI15.XI3<9>.Y XI2.XI1.XI15.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<9>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<8>.MM_i_0 VSS! XI2.XI1.XI15.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<8>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<8>.MM_i_0_15 VSS! REG_DATA_0<8> XI2.XI1.XI15.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<8>.MM_i_0_15_63 XI2.XI1.XI15.XI3<8>.DUMMY1 REG_DATA_0<8>
+ XI2.XI1.XI15.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<8>.NEN
+ XI2.XI1.XI15.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<8>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<8>.MM_i_24 VDD! XI2.XI1.XI15.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<8>.MM_i_24_1 XI2.XI1.XI15.XI3<8>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<8>.MM_i_24_0 VDD! REG_DATA_0<8> XI2.XI1.XI15.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_0<8> XI2.XI1.XI15.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI15.XI3<8>.MM_i_24_1_48 XI2.XI1.XI15.XI3<8>.Y XI2.XI1.XI15.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI15.XI3<8>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<15>.MM_i_0 VSS! XI2.XI1.XI15.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<15>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<15>.MM_i_0_15 VSS! REG_DATA_0<15> XI2.XI1.XI15.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<15>.MM_i_0_15_63 XI2.XI1.XI15.XI3<15>.DUMMY1 REG_DATA_0<15>
+ XI2.XI1.XI15.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<15>.NEN
+ XI2.XI1.XI15.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<15>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<15>.MM_i_24 VDD! XI2.XI1.XI15.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<15>.MM_i_24_1 XI2.XI1.XI15.XI3<15>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<15>.MM_i_24_0 VDD! REG_DATA_0<15> XI2.XI1.XI15.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_0<15> XI2.XI1.XI15.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<15>.MM_i_24_1_48 XI2.XI1.XI15.XI3<15>.Y
+ XI2.XI1.XI15.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI15.XI3<15>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<14>.MM_i_0 VSS! XI2.XI1.XI15.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<14>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<14>.MM_i_0_15 VSS! REG_DATA_0<14> XI2.XI1.XI15.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<14>.MM_i_0_15_63 XI2.XI1.XI15.XI3<14>.DUMMY1 REG_DATA_0<14>
+ XI2.XI1.XI15.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<14>.NEN
+ XI2.XI1.XI15.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<14>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<14>.MM_i_24 VDD! XI2.XI1.XI15.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<14>.MM_i_24_1 XI2.XI1.XI15.XI3<14>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<14>.MM_i_24_0 VDD! REG_DATA_0<14> XI2.XI1.XI15.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_0<14> XI2.XI1.XI15.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<14>.MM_i_24_1_48 XI2.XI1.XI15.XI3<14>.Y
+ XI2.XI1.XI15.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI15.XI3<14>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<13>.MM_i_0 VSS! XI2.XI1.XI15.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<13>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<13>.MM_i_0_15 VSS! REG_DATA_0<13> XI2.XI1.XI15.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<13>.MM_i_0_15_63 XI2.XI1.XI15.XI3<13>.DUMMY1 REG_DATA_0<13>
+ XI2.XI1.XI15.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<13>.NEN
+ XI2.XI1.XI15.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<13>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<13>.MM_i_24 VDD! XI2.XI1.XI15.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<13>.MM_i_24_1 XI2.XI1.XI15.XI3<13>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<13>.MM_i_24_0 VDD! REG_DATA_0<13> XI2.XI1.XI15.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_0<13> XI2.XI1.XI15.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<13>.MM_i_24_1_48 XI2.XI1.XI15.XI3<13>.Y
+ XI2.XI1.XI15.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI15.XI3<13>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI15.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI15.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI15.XI3<12>.MM_i_0 VSS! XI2.XI1.XI15.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI15.XI3<12>.MM_i_0_14 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<12>.MM_i_0_15 VSS! REG_DATA_0<12> XI2.XI1.XI15.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<12>.MM_i_0_15_63 XI2.XI1.XI15.XI3<12>.DUMMY1 REG_DATA_0<12>
+ XI2.XI1.XI15.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI15.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI15.XI3<12>.NEN
+ XI2.XI1.XI15.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI15.XI3<12>.MM_i_17 VSS! XI2.NET1<12> XI2.XI1.XI15.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI15.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI15.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<12>.MM_i_24 VDD! XI2.XI1.XI15.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI15.XI3<12>.MM_i_24_1 XI2.XI1.XI15.XI3<12>.DUMMY0 XI2.NET1<12>
+ XI2.XI1.XI15.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI15.XI3<12>.MM_i_24_0 VDD! REG_DATA_0<12> XI2.XI1.XI15.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_0<12> XI2.XI1.XI15.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI15.XI3<12>.MM_i_24_1_48 XI2.XI1.XI15.XI3<12>.Y
+ XI2.XI1.XI15.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI15.XI3<12>.MM_i_42 VDD! XI2.NET1<12> XI2.XI1.XI15.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<3>.MM_i_0 VSS! XI2.XI1.XI3.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<3>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<3>.MM_i_0_15 VSS! REG_DATA_12<3> XI2.XI1.XI3.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<3>.MM_i_0_15_63 XI2.XI1.XI3.XI3<3>.DUMMY1 REG_DATA_12<3>
+ XI2.XI1.XI3.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<3>.NEN
+ XI2.XI1.XI3.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<3>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<3>.MM_i_24 VDD! XI2.XI1.XI3.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<3>.MM_i_24_1 XI2.XI1.XI3.XI3<3>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<3>.MM_i_24_0 VDD! REG_DATA_12<3> XI2.XI1.XI3.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_12<3> XI2.XI1.XI3.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<3>.MM_i_24_1_48 XI2.XI1.XI3.XI3<3>.Y XI2.XI1.XI3.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<3>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<2>.MM_i_0 VSS! XI2.XI1.XI3.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<2>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<2>.MM_i_0_15 VSS! REG_DATA_12<2> XI2.XI1.XI3.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<2>.MM_i_0_15_63 XI2.XI1.XI3.XI3<2>.DUMMY1 REG_DATA_12<2>
+ XI2.XI1.XI3.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<2>.NEN
+ XI2.XI1.XI3.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<2>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<2>.MM_i_24 VDD! XI2.XI1.XI3.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<2>.MM_i_24_1 XI2.XI1.XI3.XI3<2>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<2>.MM_i_24_0 VDD! REG_DATA_12<2> XI2.XI1.XI3.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_12<2> XI2.XI1.XI3.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<2>.MM_i_24_1_48 XI2.XI1.XI3.XI3<2>.Y XI2.XI1.XI3.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<2>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<1>.MM_i_0 VSS! XI2.XI1.XI3.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<1>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<1>.MM_i_0_15 VSS! REG_DATA_12<1> XI2.XI1.XI3.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<1>.MM_i_0_15_63 XI2.XI1.XI3.XI3<1>.DUMMY1 REG_DATA_12<1>
+ XI2.XI1.XI3.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<1>.NEN
+ XI2.XI1.XI3.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<1>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<1>.MM_i_24 VDD! XI2.XI1.XI3.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<1>.MM_i_24_1 XI2.XI1.XI3.XI3<1>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<1>.MM_i_24_0 VDD! REG_DATA_12<1> XI2.XI1.XI3.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_12<1> XI2.XI1.XI3.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<1>.MM_i_24_1_48 XI2.XI1.XI3.XI3<1>.Y XI2.XI1.XI3.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<1>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<0>.MM_i_0 VSS! XI2.XI1.XI3.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<0>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<0>.MM_i_0_15 VSS! REG_DATA_12<0> XI2.XI1.XI3.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<0>.MM_i_0_15_63 XI2.XI1.XI3.XI3<0>.DUMMY1 REG_DATA_12<0>
+ XI2.XI1.XI3.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<0>.NEN
+ XI2.XI1.XI3.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<0>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<0>.MM_i_24 VDD! XI2.XI1.XI3.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<0>.MM_i_24_1 XI2.XI1.XI3.XI3<0>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<0>.MM_i_24_0 VDD! REG_DATA_12<0> XI2.XI1.XI3.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_12<0> XI2.XI1.XI3.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<0>.MM_i_24_1_48 XI2.XI1.XI3.XI3<0>.Y XI2.XI1.XI3.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<0>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<7>.MM_i_0 VSS! XI2.XI1.XI3.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<7>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<7>.MM_i_0_15 VSS! REG_DATA_12<7> XI2.XI1.XI3.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<7>.MM_i_0_15_63 XI2.XI1.XI3.XI3<7>.DUMMY1 REG_DATA_12<7>
+ XI2.XI1.XI3.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<7>.NEN
+ XI2.XI1.XI3.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<7>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<7>.MM_i_24 VDD! XI2.XI1.XI3.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<7>.MM_i_24_1 XI2.XI1.XI3.XI3<7>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<7>.MM_i_24_0 VDD! REG_DATA_12<7> XI2.XI1.XI3.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_12<7> XI2.XI1.XI3.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<7>.MM_i_24_1_48 XI2.XI1.XI3.XI3<7>.Y XI2.XI1.XI3.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<7>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<6>.MM_i_0 VSS! XI2.XI1.XI3.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<6>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<6>.MM_i_0_15 VSS! REG_DATA_12<6> XI2.XI1.XI3.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<6>.MM_i_0_15_63 XI2.XI1.XI3.XI3<6>.DUMMY1 REG_DATA_12<6>
+ XI2.XI1.XI3.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<6>.NEN
+ XI2.XI1.XI3.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<6>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<6>.MM_i_24 VDD! XI2.XI1.XI3.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<6>.MM_i_24_1 XI2.XI1.XI3.XI3<6>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<6>.MM_i_24_0 VDD! REG_DATA_12<6> XI2.XI1.XI3.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_12<6> XI2.XI1.XI3.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<6>.MM_i_24_1_48 XI2.XI1.XI3.XI3<6>.Y XI2.XI1.XI3.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<6>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<5>.MM_i_0 VSS! XI2.XI1.XI3.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<5>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<5>.MM_i_0_15 VSS! REG_DATA_12<5> XI2.XI1.XI3.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<5>.MM_i_0_15_63 XI2.XI1.XI3.XI3<5>.DUMMY1 REG_DATA_12<5>
+ XI2.XI1.XI3.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<5>.NEN
+ XI2.XI1.XI3.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<5>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<5>.MM_i_24 VDD! XI2.XI1.XI3.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<5>.MM_i_24_1 XI2.XI1.XI3.XI3<5>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<5>.MM_i_24_0 VDD! REG_DATA_12<5> XI2.XI1.XI3.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_12<5> XI2.XI1.XI3.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<5>.MM_i_24_1_48 XI2.XI1.XI3.XI3<5>.Y XI2.XI1.XI3.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<5>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<4>.MM_i_0 VSS! XI2.XI1.XI3.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<4>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<4>.MM_i_0_15 VSS! REG_DATA_12<4> XI2.XI1.XI3.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<4>.MM_i_0_15_63 XI2.XI1.XI3.XI3<4>.DUMMY1 REG_DATA_12<4>
+ XI2.XI1.XI3.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<4>.NEN
+ XI2.XI1.XI3.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<4>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<4>.MM_i_24 VDD! XI2.XI1.XI3.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<4>.MM_i_24_1 XI2.XI1.XI3.XI3<4>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<4>.MM_i_24_0 VDD! REG_DATA_12<4> XI2.XI1.XI3.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_12<4> XI2.XI1.XI3.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<4>.MM_i_24_1_48 XI2.XI1.XI3.XI3<4>.Y XI2.XI1.XI3.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<4>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<11>.MM_i_0 VSS! XI2.XI1.XI3.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<11>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<11>.MM_i_0_15 VSS! REG_DATA_12<11> XI2.XI1.XI3.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<11>.MM_i_0_15_63 XI2.XI1.XI3.XI3<11>.DUMMY1 REG_DATA_12<11>
+ XI2.XI1.XI3.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<11>.NEN
+ XI2.XI1.XI3.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<11>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<11>.MM_i_24 VDD! XI2.XI1.XI3.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<11>.MM_i_24_1 XI2.XI1.XI3.XI3<11>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<11>.MM_i_24_0 VDD! REG_DATA_12<11> XI2.XI1.XI3.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_12<11> XI2.XI1.XI3.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<11>.MM_i_24_1_48 XI2.XI1.XI3.XI3<11>.Y XI2.XI1.XI3.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<11>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<10>.MM_i_0 VSS! XI2.XI1.XI3.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<10>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<10>.MM_i_0_15 VSS! REG_DATA_12<10> XI2.XI1.XI3.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<10>.MM_i_0_15_63 XI2.XI1.XI3.XI3<10>.DUMMY1 REG_DATA_12<10>
+ XI2.XI1.XI3.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<10>.NEN
+ XI2.XI1.XI3.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<10>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<10>.MM_i_24 VDD! XI2.XI1.XI3.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<10>.MM_i_24_1 XI2.XI1.XI3.XI3<10>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<10>.MM_i_24_0 VDD! REG_DATA_12<10> XI2.XI1.XI3.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_12<10> XI2.XI1.XI3.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<10>.MM_i_24_1_48 XI2.XI1.XI3.XI3<10>.Y XI2.XI1.XI3.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<10>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<9>.MM_i_0 VSS! XI2.XI1.XI3.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<9>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<9>.MM_i_0_15 VSS! REG_DATA_12<9> XI2.XI1.XI3.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<9>.MM_i_0_15_63 XI2.XI1.XI3.XI3<9>.DUMMY1 REG_DATA_12<9>
+ XI2.XI1.XI3.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<9>.NEN
+ XI2.XI1.XI3.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<9>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<9>.MM_i_24 VDD! XI2.XI1.XI3.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<9>.MM_i_24_1 XI2.XI1.XI3.XI3<9>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<9>.MM_i_24_0 VDD! REG_DATA_12<9> XI2.XI1.XI3.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_12<9> XI2.XI1.XI3.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<9>.MM_i_24_1_48 XI2.XI1.XI3.XI3<9>.Y XI2.XI1.XI3.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<9>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<8>.MM_i_0 VSS! XI2.XI1.XI3.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<8>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<8>.MM_i_0_15 VSS! REG_DATA_12<8> XI2.XI1.XI3.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<8>.MM_i_0_15_63 XI2.XI1.XI3.XI3<8>.DUMMY1 REG_DATA_12<8>
+ XI2.XI1.XI3.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<8>.NEN
+ XI2.XI1.XI3.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<8>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<8>.MM_i_24 VDD! XI2.XI1.XI3.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<8>.MM_i_24_1 XI2.XI1.XI3.XI3<8>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<8>.MM_i_24_0 VDD! REG_DATA_12<8> XI2.XI1.XI3.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_12<8> XI2.XI1.XI3.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI3.XI3<8>.MM_i_24_1_48 XI2.XI1.XI3.XI3<8>.Y XI2.XI1.XI3.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<8>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<15>.MM_i_0 VSS! XI2.XI1.XI3.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<15>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<15>.MM_i_0_15 VSS! REG_DATA_12<15> XI2.XI1.XI3.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<15>.MM_i_0_15_63 XI2.XI1.XI3.XI3<15>.DUMMY1 REG_DATA_12<15>
+ XI2.XI1.XI3.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<15>.NEN
+ XI2.XI1.XI3.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<15>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<15>.MM_i_24 VDD! XI2.XI1.XI3.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<15>.MM_i_24_1 XI2.XI1.XI3.XI3<15>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<15>.MM_i_24_0 VDD! REG_DATA_12<15> XI2.XI1.XI3.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_12<15> XI2.XI1.XI3.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<15>.MM_i_24_1_48 XI2.XI1.XI3.XI3<15>.Y XI2.XI1.XI3.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<15>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<14>.MM_i_0 VSS! XI2.XI1.XI3.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<14>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<14>.MM_i_0_15 VSS! REG_DATA_12<14> XI2.XI1.XI3.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<14>.MM_i_0_15_63 XI2.XI1.XI3.XI3<14>.DUMMY1 REG_DATA_12<14>
+ XI2.XI1.XI3.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<14>.NEN
+ XI2.XI1.XI3.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<14>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<14>.MM_i_24 VDD! XI2.XI1.XI3.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<14>.MM_i_24_1 XI2.XI1.XI3.XI3<14>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<14>.MM_i_24_0 VDD! REG_DATA_12<14> XI2.XI1.XI3.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_12<14> XI2.XI1.XI3.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<14>.MM_i_24_1_48 XI2.XI1.XI3.XI3<14>.Y XI2.XI1.XI3.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<14>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<13>.MM_i_0 VSS! XI2.XI1.XI3.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<13>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<13>.MM_i_0_15 VSS! REG_DATA_12<13> XI2.XI1.XI3.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<13>.MM_i_0_15_63 XI2.XI1.XI3.XI3<13>.DUMMY1 REG_DATA_12<13>
+ XI2.XI1.XI3.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<13>.NEN
+ XI2.XI1.XI3.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<13>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<13>.MM_i_24 VDD! XI2.XI1.XI3.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<13>.MM_i_24_1 XI2.XI1.XI3.XI3<13>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<13>.MM_i_24_0 VDD! REG_DATA_12<13> XI2.XI1.XI3.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_12<13> XI2.XI1.XI3.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<13>.MM_i_24_1_48 XI2.XI1.XI3.XI3<13>.Y XI2.XI1.XI3.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<13>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI3.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI3.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI3.XI3<12>.MM_i_0 VSS! XI2.XI1.XI3.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI3.XI3<12>.MM_i_0_14 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<12>.MM_i_0_15 VSS! REG_DATA_12<12> XI2.XI1.XI3.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<12>.MM_i_0_15_63 XI2.XI1.XI3.XI3<12>.DUMMY1 REG_DATA_12<12>
+ XI2.XI1.XI3.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI3.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI3.XI3<12>.NEN
+ XI2.XI1.XI3.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI3.XI3<12>.MM_i_17 VSS! XI2.NET1<0> XI2.XI1.XI3.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI3.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI3.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<12>.MM_i_24 VDD! XI2.XI1.XI3.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI3.XI3<12>.MM_i_24_1 XI2.XI1.XI3.XI3<12>.DUMMY0 XI2.NET1<0>
+ XI2.XI1.XI3.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI3.XI3<12>.MM_i_24_0 VDD! REG_DATA_12<12> XI2.XI1.XI3.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_12<12> XI2.XI1.XI3.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI3.XI3<12>.MM_i_24_1_48 XI2.XI1.XI3.XI3<12>.Y XI2.XI1.XI3.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI3.XI3<12>.MM_i_42 VDD! XI2.NET1<0> XI2.XI1.XI3.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<3>.MM_i_0 VSS! XI2.XI1.XI4.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<3>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<3>.MM_i_0_15 VSS! REG_DATA_11<3> XI2.XI1.XI4.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<3>.MM_i_0_15_63 XI2.XI1.XI4.XI3<3>.DUMMY1 REG_DATA_11<3>
+ XI2.XI1.XI4.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<3>.NEN
+ XI2.XI1.XI4.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<3>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<3>.MM_i_24 VDD! XI2.XI1.XI4.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<3>.MM_i_24_1 XI2.XI1.XI4.XI3<3>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<3>.MM_i_24_0 VDD! REG_DATA_11<3> XI2.XI1.XI4.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_11<3> XI2.XI1.XI4.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<3>.MM_i_24_1_48 XI2.XI1.XI4.XI3<3>.Y XI2.XI1.XI4.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<3>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<2>.MM_i_0 VSS! XI2.XI1.XI4.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<2>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<2>.MM_i_0_15 VSS! REG_DATA_11<2> XI2.XI1.XI4.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<2>.MM_i_0_15_63 XI2.XI1.XI4.XI3<2>.DUMMY1 REG_DATA_11<2>
+ XI2.XI1.XI4.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<2>.NEN
+ XI2.XI1.XI4.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<2>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<2>.MM_i_24 VDD! XI2.XI1.XI4.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<2>.MM_i_24_1 XI2.XI1.XI4.XI3<2>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<2>.MM_i_24_0 VDD! REG_DATA_11<2> XI2.XI1.XI4.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_11<2> XI2.XI1.XI4.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<2>.MM_i_24_1_48 XI2.XI1.XI4.XI3<2>.Y XI2.XI1.XI4.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<2>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<1>.MM_i_0 VSS! XI2.XI1.XI4.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<1>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<1>.MM_i_0_15 VSS! REG_DATA_11<1> XI2.XI1.XI4.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<1>.MM_i_0_15_63 XI2.XI1.XI4.XI3<1>.DUMMY1 REG_DATA_11<1>
+ XI2.XI1.XI4.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<1>.NEN
+ XI2.XI1.XI4.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<1>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<1>.MM_i_24 VDD! XI2.XI1.XI4.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<1>.MM_i_24_1 XI2.XI1.XI4.XI3<1>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<1>.MM_i_24_0 VDD! REG_DATA_11<1> XI2.XI1.XI4.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_11<1> XI2.XI1.XI4.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<1>.MM_i_24_1_48 XI2.XI1.XI4.XI3<1>.Y XI2.XI1.XI4.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<1>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<0>.MM_i_0 VSS! XI2.XI1.XI4.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<0>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<0>.MM_i_0_15 VSS! REG_DATA_11<0> XI2.XI1.XI4.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<0>.MM_i_0_15_63 XI2.XI1.XI4.XI3<0>.DUMMY1 REG_DATA_11<0>
+ XI2.XI1.XI4.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<0>.NEN
+ XI2.XI1.XI4.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<0>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<0>.MM_i_24 VDD! XI2.XI1.XI4.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<0>.MM_i_24_1 XI2.XI1.XI4.XI3<0>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<0>.MM_i_24_0 VDD! REG_DATA_11<0> XI2.XI1.XI4.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_11<0> XI2.XI1.XI4.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<0>.MM_i_24_1_48 XI2.XI1.XI4.XI3<0>.Y XI2.XI1.XI4.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<0>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<7>.MM_i_0 VSS! XI2.XI1.XI4.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<7>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<7>.MM_i_0_15 VSS! REG_DATA_11<7> XI2.XI1.XI4.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<7>.MM_i_0_15_63 XI2.XI1.XI4.XI3<7>.DUMMY1 REG_DATA_11<7>
+ XI2.XI1.XI4.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<7>.NEN
+ XI2.XI1.XI4.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<7>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<7>.MM_i_24 VDD! XI2.XI1.XI4.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<7>.MM_i_24_1 XI2.XI1.XI4.XI3<7>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<7>.MM_i_24_0 VDD! REG_DATA_11<7> XI2.XI1.XI4.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_11<7> XI2.XI1.XI4.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<7>.MM_i_24_1_48 XI2.XI1.XI4.XI3<7>.Y XI2.XI1.XI4.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<7>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<6>.MM_i_0 VSS! XI2.XI1.XI4.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<6>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<6>.MM_i_0_15 VSS! REG_DATA_11<6> XI2.XI1.XI4.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<6>.MM_i_0_15_63 XI2.XI1.XI4.XI3<6>.DUMMY1 REG_DATA_11<6>
+ XI2.XI1.XI4.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<6>.NEN
+ XI2.XI1.XI4.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<6>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<6>.MM_i_24 VDD! XI2.XI1.XI4.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<6>.MM_i_24_1 XI2.XI1.XI4.XI3<6>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<6>.MM_i_24_0 VDD! REG_DATA_11<6> XI2.XI1.XI4.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_11<6> XI2.XI1.XI4.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<6>.MM_i_24_1_48 XI2.XI1.XI4.XI3<6>.Y XI2.XI1.XI4.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<6>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<5>.MM_i_0 VSS! XI2.XI1.XI4.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<5>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<5>.MM_i_0_15 VSS! REG_DATA_11<5> XI2.XI1.XI4.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<5>.MM_i_0_15_63 XI2.XI1.XI4.XI3<5>.DUMMY1 REG_DATA_11<5>
+ XI2.XI1.XI4.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<5>.NEN
+ XI2.XI1.XI4.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<5>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<5>.MM_i_24 VDD! XI2.XI1.XI4.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<5>.MM_i_24_1 XI2.XI1.XI4.XI3<5>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<5>.MM_i_24_0 VDD! REG_DATA_11<5> XI2.XI1.XI4.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_11<5> XI2.XI1.XI4.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<5>.MM_i_24_1_48 XI2.XI1.XI4.XI3<5>.Y XI2.XI1.XI4.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<5>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<4>.MM_i_0 VSS! XI2.XI1.XI4.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<4>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<4>.MM_i_0_15 VSS! REG_DATA_11<4> XI2.XI1.XI4.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<4>.MM_i_0_15_63 XI2.XI1.XI4.XI3<4>.DUMMY1 REG_DATA_11<4>
+ XI2.XI1.XI4.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<4>.NEN
+ XI2.XI1.XI4.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<4>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<4>.MM_i_24 VDD! XI2.XI1.XI4.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<4>.MM_i_24_1 XI2.XI1.XI4.XI3<4>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<4>.MM_i_24_0 VDD! REG_DATA_11<4> XI2.XI1.XI4.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_11<4> XI2.XI1.XI4.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<4>.MM_i_24_1_48 XI2.XI1.XI4.XI3<4>.Y XI2.XI1.XI4.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<4>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<11>.MM_i_0 VSS! XI2.XI1.XI4.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<11>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<11>.MM_i_0_15 VSS! REG_DATA_11<11> XI2.XI1.XI4.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<11>.MM_i_0_15_63 XI2.XI1.XI4.XI3<11>.DUMMY1 REG_DATA_11<11>
+ XI2.XI1.XI4.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<11>.NEN
+ XI2.XI1.XI4.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<11>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<11>.MM_i_24 VDD! XI2.XI1.XI4.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<11>.MM_i_24_1 XI2.XI1.XI4.XI3<11>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<11>.MM_i_24_0 VDD! REG_DATA_11<11> XI2.XI1.XI4.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_11<11> XI2.XI1.XI4.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<11>.MM_i_24_1_48 XI2.XI1.XI4.XI3<11>.Y XI2.XI1.XI4.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<11>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<10>.MM_i_0 VSS! XI2.XI1.XI4.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<10>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<10>.MM_i_0_15 VSS! REG_DATA_11<10> XI2.XI1.XI4.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<10>.MM_i_0_15_63 XI2.XI1.XI4.XI3<10>.DUMMY1 REG_DATA_11<10>
+ XI2.XI1.XI4.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<10>.NEN
+ XI2.XI1.XI4.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<10>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<10>.MM_i_24 VDD! XI2.XI1.XI4.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<10>.MM_i_24_1 XI2.XI1.XI4.XI3<10>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<10>.MM_i_24_0 VDD! REG_DATA_11<10> XI2.XI1.XI4.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_11<10> XI2.XI1.XI4.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<10>.MM_i_24_1_48 XI2.XI1.XI4.XI3<10>.Y XI2.XI1.XI4.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<10>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<9>.MM_i_0 VSS! XI2.XI1.XI4.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<9>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<9>.MM_i_0_15 VSS! REG_DATA_11<9> XI2.XI1.XI4.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<9>.MM_i_0_15_63 XI2.XI1.XI4.XI3<9>.DUMMY1 REG_DATA_11<9>
+ XI2.XI1.XI4.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<9>.NEN
+ XI2.XI1.XI4.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<9>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<9>.MM_i_24 VDD! XI2.XI1.XI4.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<9>.MM_i_24_1 XI2.XI1.XI4.XI3<9>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<9>.MM_i_24_0 VDD! REG_DATA_11<9> XI2.XI1.XI4.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_11<9> XI2.XI1.XI4.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<9>.MM_i_24_1_48 XI2.XI1.XI4.XI3<9>.Y XI2.XI1.XI4.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<9>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<8>.MM_i_0 VSS! XI2.XI1.XI4.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<8>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<8>.MM_i_0_15 VSS! REG_DATA_11<8> XI2.XI1.XI4.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<8>.MM_i_0_15_63 XI2.XI1.XI4.XI3<8>.DUMMY1 REG_DATA_11<8>
+ XI2.XI1.XI4.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<8>.NEN
+ XI2.XI1.XI4.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<8>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<8>.MM_i_24 VDD! XI2.XI1.XI4.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<8>.MM_i_24_1 XI2.XI1.XI4.XI3<8>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<8>.MM_i_24_0 VDD! REG_DATA_11<8> XI2.XI1.XI4.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_11<8> XI2.XI1.XI4.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI4.XI3<8>.MM_i_24_1_48 XI2.XI1.XI4.XI3<8>.Y XI2.XI1.XI4.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<8>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<15>.MM_i_0 VSS! XI2.XI1.XI4.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<15>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<15>.MM_i_0_15 VSS! REG_DATA_11<15> XI2.XI1.XI4.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<15>.MM_i_0_15_63 XI2.XI1.XI4.XI3<15>.DUMMY1 REG_DATA_11<15>
+ XI2.XI1.XI4.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<15>.NEN
+ XI2.XI1.XI4.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<15>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<15>.MM_i_24 VDD! XI2.XI1.XI4.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<15>.MM_i_24_1 XI2.XI1.XI4.XI3<15>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<15>.MM_i_24_0 VDD! REG_DATA_11<15> XI2.XI1.XI4.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_11<15> XI2.XI1.XI4.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<15>.MM_i_24_1_48 XI2.XI1.XI4.XI3<15>.Y XI2.XI1.XI4.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<15>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<14>.MM_i_0 VSS! XI2.XI1.XI4.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<14>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<14>.MM_i_0_15 VSS! REG_DATA_11<14> XI2.XI1.XI4.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<14>.MM_i_0_15_63 XI2.XI1.XI4.XI3<14>.DUMMY1 REG_DATA_11<14>
+ XI2.XI1.XI4.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<14>.NEN
+ XI2.XI1.XI4.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<14>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<14>.MM_i_24 VDD! XI2.XI1.XI4.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<14>.MM_i_24_1 XI2.XI1.XI4.XI3<14>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<14>.MM_i_24_0 VDD! REG_DATA_11<14> XI2.XI1.XI4.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_11<14> XI2.XI1.XI4.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<14>.MM_i_24_1_48 XI2.XI1.XI4.XI3<14>.Y XI2.XI1.XI4.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<14>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<13>.MM_i_0 VSS! XI2.XI1.XI4.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<13>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<13>.MM_i_0_15 VSS! REG_DATA_11<13> XI2.XI1.XI4.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<13>.MM_i_0_15_63 XI2.XI1.XI4.XI3<13>.DUMMY1 REG_DATA_11<13>
+ XI2.XI1.XI4.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<13>.NEN
+ XI2.XI1.XI4.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<13>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<13>.MM_i_24 VDD! XI2.XI1.XI4.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<13>.MM_i_24_1 XI2.XI1.XI4.XI3<13>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<13>.MM_i_24_0 VDD! REG_DATA_11<13> XI2.XI1.XI4.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_11<13> XI2.XI1.XI4.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<13>.MM_i_24_1_48 XI2.XI1.XI4.XI3<13>.Y XI2.XI1.XI4.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<13>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI4.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI4.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI4.XI3<12>.MM_i_0 VSS! XI2.XI1.XI4.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI4.XI3<12>.MM_i_0_14 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<12>.MM_i_0_15 VSS! REG_DATA_11<12> XI2.XI1.XI4.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<12>.MM_i_0_15_63 XI2.XI1.XI4.XI3<12>.DUMMY1 REG_DATA_11<12>
+ XI2.XI1.XI4.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI4.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI4.XI3<12>.NEN
+ XI2.XI1.XI4.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI4.XI3<12>.MM_i_17 VSS! XI2.NET1<1> XI2.XI1.XI4.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI4.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI4.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<12>.MM_i_24 VDD! XI2.XI1.XI4.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI4.XI3<12>.MM_i_24_1 XI2.XI1.XI4.XI3<12>.DUMMY0 XI2.NET1<1>
+ XI2.XI1.XI4.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI4.XI3<12>.MM_i_24_0 VDD! REG_DATA_11<12> XI2.XI1.XI4.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_11<12> XI2.XI1.XI4.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI4.XI3<12>.MM_i_24_1_48 XI2.XI1.XI4.XI3<12>.Y XI2.XI1.XI4.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI4.XI3<12>.MM_i_42 VDD! XI2.NET1<1> XI2.XI1.XI4.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<3>.MM_i_0 VSS! XI2.XI1.XI6.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<3>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<3>.MM_i_0_15 VSS! REG_DATA_10<3> XI2.XI1.XI6.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<3>.MM_i_0_15_63 XI2.XI1.XI6.XI3<3>.DUMMY1 REG_DATA_10<3>
+ XI2.XI1.XI6.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<3>.NEN
+ XI2.XI1.XI6.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<3>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<3>.MM_i_24 VDD! XI2.XI1.XI6.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<3>.MM_i_24_1 XI2.XI1.XI6.XI3<3>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<3>.MM_i_24_0 VDD! REG_DATA_10<3> XI2.XI1.XI6.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_10<3> XI2.XI1.XI6.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<3>.MM_i_24_1_48 XI2.XI1.XI6.XI3<3>.Y XI2.XI1.XI6.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<3>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<2>.MM_i_0 VSS! XI2.XI1.XI6.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<2>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<2>.MM_i_0_15 VSS! REG_DATA_10<2> XI2.XI1.XI6.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<2>.MM_i_0_15_63 XI2.XI1.XI6.XI3<2>.DUMMY1 REG_DATA_10<2>
+ XI2.XI1.XI6.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<2>.NEN
+ XI2.XI1.XI6.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<2>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<2>.MM_i_24 VDD! XI2.XI1.XI6.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<2>.MM_i_24_1 XI2.XI1.XI6.XI3<2>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<2>.MM_i_24_0 VDD! REG_DATA_10<2> XI2.XI1.XI6.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_10<2> XI2.XI1.XI6.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<2>.MM_i_24_1_48 XI2.XI1.XI6.XI3<2>.Y XI2.XI1.XI6.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<2>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<1>.MM_i_0 VSS! XI2.XI1.XI6.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<1>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<1>.MM_i_0_15 VSS! REG_DATA_10<1> XI2.XI1.XI6.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<1>.MM_i_0_15_63 XI2.XI1.XI6.XI3<1>.DUMMY1 REG_DATA_10<1>
+ XI2.XI1.XI6.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<1>.NEN
+ XI2.XI1.XI6.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<1>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<1>.MM_i_24 VDD! XI2.XI1.XI6.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<1>.MM_i_24_1 XI2.XI1.XI6.XI3<1>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<1>.MM_i_24_0 VDD! REG_DATA_10<1> XI2.XI1.XI6.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_10<1> XI2.XI1.XI6.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<1>.MM_i_24_1_48 XI2.XI1.XI6.XI3<1>.Y XI2.XI1.XI6.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<1>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<0>.MM_i_0 VSS! XI2.XI1.XI6.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<0>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<0>.MM_i_0_15 VSS! REG_DATA_10<0> XI2.XI1.XI6.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<0>.MM_i_0_15_63 XI2.XI1.XI6.XI3<0>.DUMMY1 REG_DATA_10<0>
+ XI2.XI1.XI6.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<0>.NEN
+ XI2.XI1.XI6.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<0>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<0>.MM_i_24 VDD! XI2.XI1.XI6.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<0>.MM_i_24_1 XI2.XI1.XI6.XI3<0>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<0>.MM_i_24_0 VDD! REG_DATA_10<0> XI2.XI1.XI6.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_10<0> XI2.XI1.XI6.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<0>.MM_i_24_1_48 XI2.XI1.XI6.XI3<0>.Y XI2.XI1.XI6.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<0>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<7>.MM_i_0 VSS! XI2.XI1.XI6.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<7>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<7>.MM_i_0_15 VSS! REG_DATA_10<7> XI2.XI1.XI6.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<7>.MM_i_0_15_63 XI2.XI1.XI6.XI3<7>.DUMMY1 REG_DATA_10<7>
+ XI2.XI1.XI6.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<7>.NEN
+ XI2.XI1.XI6.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<7>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<7>.MM_i_24 VDD! XI2.XI1.XI6.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<7>.MM_i_24_1 XI2.XI1.XI6.XI3<7>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<7>.MM_i_24_0 VDD! REG_DATA_10<7> XI2.XI1.XI6.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_10<7> XI2.XI1.XI6.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<7>.MM_i_24_1_48 XI2.XI1.XI6.XI3<7>.Y XI2.XI1.XI6.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<7>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<6>.MM_i_0 VSS! XI2.XI1.XI6.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<6>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<6>.MM_i_0_15 VSS! REG_DATA_10<6> XI2.XI1.XI6.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<6>.MM_i_0_15_63 XI2.XI1.XI6.XI3<6>.DUMMY1 REG_DATA_10<6>
+ XI2.XI1.XI6.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<6>.NEN
+ XI2.XI1.XI6.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<6>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<6>.MM_i_24 VDD! XI2.XI1.XI6.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<6>.MM_i_24_1 XI2.XI1.XI6.XI3<6>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<6>.MM_i_24_0 VDD! REG_DATA_10<6> XI2.XI1.XI6.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_10<6> XI2.XI1.XI6.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<6>.MM_i_24_1_48 XI2.XI1.XI6.XI3<6>.Y XI2.XI1.XI6.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<6>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<5>.MM_i_0 VSS! XI2.XI1.XI6.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<5>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<5>.MM_i_0_15 VSS! REG_DATA_10<5> XI2.XI1.XI6.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<5>.MM_i_0_15_63 XI2.XI1.XI6.XI3<5>.DUMMY1 REG_DATA_10<5>
+ XI2.XI1.XI6.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<5>.NEN
+ XI2.XI1.XI6.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<5>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<5>.MM_i_24 VDD! XI2.XI1.XI6.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<5>.MM_i_24_1 XI2.XI1.XI6.XI3<5>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<5>.MM_i_24_0 VDD! REG_DATA_10<5> XI2.XI1.XI6.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_10<5> XI2.XI1.XI6.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<5>.MM_i_24_1_48 XI2.XI1.XI6.XI3<5>.Y XI2.XI1.XI6.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<5>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<4>.MM_i_0 VSS! XI2.XI1.XI6.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<4>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<4>.MM_i_0_15 VSS! REG_DATA_10<4> XI2.XI1.XI6.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<4>.MM_i_0_15_63 XI2.XI1.XI6.XI3<4>.DUMMY1 REG_DATA_10<4>
+ XI2.XI1.XI6.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<4>.NEN
+ XI2.XI1.XI6.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<4>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<4>.MM_i_24 VDD! XI2.XI1.XI6.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<4>.MM_i_24_1 XI2.XI1.XI6.XI3<4>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<4>.MM_i_24_0 VDD! REG_DATA_10<4> XI2.XI1.XI6.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_10<4> XI2.XI1.XI6.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<4>.MM_i_24_1_48 XI2.XI1.XI6.XI3<4>.Y XI2.XI1.XI6.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<4>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<11>.MM_i_0 VSS! XI2.XI1.XI6.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<11>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<11>.MM_i_0_15 VSS! REG_DATA_10<11> XI2.XI1.XI6.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<11>.MM_i_0_15_63 XI2.XI1.XI6.XI3<11>.DUMMY1 REG_DATA_10<11>
+ XI2.XI1.XI6.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<11>.NEN
+ XI2.XI1.XI6.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<11>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<11>.MM_i_24 VDD! XI2.XI1.XI6.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<11>.MM_i_24_1 XI2.XI1.XI6.XI3<11>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<11>.MM_i_24_0 VDD! REG_DATA_10<11> XI2.XI1.XI6.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_10<11> XI2.XI1.XI6.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<11>.MM_i_24_1_48 XI2.XI1.XI6.XI3<11>.Y XI2.XI1.XI6.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<11>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<10>.MM_i_0 VSS! XI2.XI1.XI6.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<10>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<10>.MM_i_0_15 VSS! REG_DATA_10<10> XI2.XI1.XI6.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<10>.MM_i_0_15_63 XI2.XI1.XI6.XI3<10>.DUMMY1 REG_DATA_10<10>
+ XI2.XI1.XI6.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<10>.NEN
+ XI2.XI1.XI6.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<10>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<10>.MM_i_24 VDD! XI2.XI1.XI6.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<10>.MM_i_24_1 XI2.XI1.XI6.XI3<10>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<10>.MM_i_24_0 VDD! REG_DATA_10<10> XI2.XI1.XI6.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_10<10> XI2.XI1.XI6.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<10>.MM_i_24_1_48 XI2.XI1.XI6.XI3<10>.Y XI2.XI1.XI6.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<10>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<9>.MM_i_0 VSS! XI2.XI1.XI6.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<9>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<9>.MM_i_0_15 VSS! REG_DATA_10<9> XI2.XI1.XI6.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<9>.MM_i_0_15_63 XI2.XI1.XI6.XI3<9>.DUMMY1 REG_DATA_10<9>
+ XI2.XI1.XI6.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<9>.NEN
+ XI2.XI1.XI6.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<9>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<9>.MM_i_24 VDD! XI2.XI1.XI6.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<9>.MM_i_24_1 XI2.XI1.XI6.XI3<9>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<9>.MM_i_24_0 VDD! REG_DATA_10<9> XI2.XI1.XI6.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_10<9> XI2.XI1.XI6.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<9>.MM_i_24_1_48 XI2.XI1.XI6.XI3<9>.Y XI2.XI1.XI6.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<9>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<8>.MM_i_0 VSS! XI2.XI1.XI6.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<8>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<8>.MM_i_0_15 VSS! REG_DATA_10<8> XI2.XI1.XI6.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<8>.MM_i_0_15_63 XI2.XI1.XI6.XI3<8>.DUMMY1 REG_DATA_10<8>
+ XI2.XI1.XI6.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<8>.NEN
+ XI2.XI1.XI6.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<8>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<8>.MM_i_24 VDD! XI2.XI1.XI6.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<8>.MM_i_24_1 XI2.XI1.XI6.XI3<8>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<8>.MM_i_24_0 VDD! REG_DATA_10<8> XI2.XI1.XI6.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_10<8> XI2.XI1.XI6.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI6.XI3<8>.MM_i_24_1_48 XI2.XI1.XI6.XI3<8>.Y XI2.XI1.XI6.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<8>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<15>.MM_i_0 VSS! XI2.XI1.XI6.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<15>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<15>.MM_i_0_15 VSS! REG_DATA_10<15> XI2.XI1.XI6.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<15>.MM_i_0_15_63 XI2.XI1.XI6.XI3<15>.DUMMY1 REG_DATA_10<15>
+ XI2.XI1.XI6.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<15>.NEN
+ XI2.XI1.XI6.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<15>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<15>.MM_i_24 VDD! XI2.XI1.XI6.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<15>.MM_i_24_1 XI2.XI1.XI6.XI3<15>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<15>.MM_i_24_0 VDD! REG_DATA_10<15> XI2.XI1.XI6.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_10<15> XI2.XI1.XI6.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<15>.MM_i_24_1_48 XI2.XI1.XI6.XI3<15>.Y XI2.XI1.XI6.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<15>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<14>.MM_i_0 VSS! XI2.XI1.XI6.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<14>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<14>.MM_i_0_15 VSS! REG_DATA_10<14> XI2.XI1.XI6.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<14>.MM_i_0_15_63 XI2.XI1.XI6.XI3<14>.DUMMY1 REG_DATA_10<14>
+ XI2.XI1.XI6.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<14>.NEN
+ XI2.XI1.XI6.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<14>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<14>.MM_i_24 VDD! XI2.XI1.XI6.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<14>.MM_i_24_1 XI2.XI1.XI6.XI3<14>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<14>.MM_i_24_0 VDD! REG_DATA_10<14> XI2.XI1.XI6.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_10<14> XI2.XI1.XI6.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<14>.MM_i_24_1_48 XI2.XI1.XI6.XI3<14>.Y XI2.XI1.XI6.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<14>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<13>.MM_i_0 VSS! XI2.XI1.XI6.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<13>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<13>.MM_i_0_15 VSS! REG_DATA_10<13> XI2.XI1.XI6.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<13>.MM_i_0_15_63 XI2.XI1.XI6.XI3<13>.DUMMY1 REG_DATA_10<13>
+ XI2.XI1.XI6.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<13>.NEN
+ XI2.XI1.XI6.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<13>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<13>.MM_i_24 VDD! XI2.XI1.XI6.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<13>.MM_i_24_1 XI2.XI1.XI6.XI3<13>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<13>.MM_i_24_0 VDD! REG_DATA_10<13> XI2.XI1.XI6.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_10<13> XI2.XI1.XI6.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<13>.MM_i_24_1_48 XI2.XI1.XI6.XI3<13>.Y XI2.XI1.XI6.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<13>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI6.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI6.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI6.XI3<12>.MM_i_0 VSS! XI2.XI1.XI6.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI6.XI3<12>.MM_i_0_14 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<12>.MM_i_0_15 VSS! REG_DATA_10<12> XI2.XI1.XI6.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<12>.MM_i_0_15_63 XI2.XI1.XI6.XI3<12>.DUMMY1 REG_DATA_10<12>
+ XI2.XI1.XI6.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI6.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI6.XI3<12>.NEN
+ XI2.XI1.XI6.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI6.XI3<12>.MM_i_17 VSS! XI2.NET1<2> XI2.XI1.XI6.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI6.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI6.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<12>.MM_i_24 VDD! XI2.XI1.XI6.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI6.XI3<12>.MM_i_24_1 XI2.XI1.XI6.XI3<12>.DUMMY0 XI2.NET1<2>
+ XI2.XI1.XI6.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI6.XI3<12>.MM_i_24_0 VDD! REG_DATA_10<12> XI2.XI1.XI6.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_10<12> XI2.XI1.XI6.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI6.XI3<12>.MM_i_24_1_48 XI2.XI1.XI6.XI3<12>.Y XI2.XI1.XI6.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI6.XI3<12>.MM_i_42 VDD! XI2.NET1<2> XI2.XI1.XI6.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<3>.MM_i_0 VSS! XI2.XI1.XI5.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<3>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<3>.MM_i_0_15 VSS! REG_DATA_9<3> XI2.XI1.XI5.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<3>.MM_i_0_15_63 XI2.XI1.XI5.XI3<3>.DUMMY1 REG_DATA_9<3>
+ XI2.XI1.XI5.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<3>.NEN
+ XI2.XI1.XI5.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<3>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<3>.MM_i_24 VDD! XI2.XI1.XI5.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<3>.MM_i_24_1 XI2.XI1.XI5.XI3<3>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<3>.MM_i_24_0 VDD! REG_DATA_9<3> XI2.XI1.XI5.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_9<3> XI2.XI1.XI5.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<3>.MM_i_24_1_48 XI2.XI1.XI5.XI3<3>.Y XI2.XI1.XI5.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<3>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<2>.MM_i_0 VSS! XI2.XI1.XI5.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<2>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<2>.MM_i_0_15 VSS! REG_DATA_9<2> XI2.XI1.XI5.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<2>.MM_i_0_15_63 XI2.XI1.XI5.XI3<2>.DUMMY1 REG_DATA_9<2>
+ XI2.XI1.XI5.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<2>.NEN
+ XI2.XI1.XI5.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<2>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<2>.MM_i_24 VDD! XI2.XI1.XI5.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<2>.MM_i_24_1 XI2.XI1.XI5.XI3<2>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<2>.MM_i_24_0 VDD! REG_DATA_9<2> XI2.XI1.XI5.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_9<2> XI2.XI1.XI5.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<2>.MM_i_24_1_48 XI2.XI1.XI5.XI3<2>.Y XI2.XI1.XI5.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<2>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<1>.MM_i_0 VSS! XI2.XI1.XI5.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<1>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<1>.MM_i_0_15 VSS! REG_DATA_9<1> XI2.XI1.XI5.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<1>.MM_i_0_15_63 XI2.XI1.XI5.XI3<1>.DUMMY1 REG_DATA_9<1>
+ XI2.XI1.XI5.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<1>.NEN
+ XI2.XI1.XI5.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<1>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<1>.MM_i_24 VDD! XI2.XI1.XI5.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<1>.MM_i_24_1 XI2.XI1.XI5.XI3<1>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<1>.MM_i_24_0 VDD! REG_DATA_9<1> XI2.XI1.XI5.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_9<1> XI2.XI1.XI5.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<1>.MM_i_24_1_48 XI2.XI1.XI5.XI3<1>.Y XI2.XI1.XI5.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<1>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<0>.MM_i_0 VSS! XI2.XI1.XI5.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<0>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<0>.MM_i_0_15 VSS! REG_DATA_9<0> XI2.XI1.XI5.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<0>.MM_i_0_15_63 XI2.XI1.XI5.XI3<0>.DUMMY1 REG_DATA_9<0>
+ XI2.XI1.XI5.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<0>.NEN
+ XI2.XI1.XI5.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<0>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<0>.MM_i_24 VDD! XI2.XI1.XI5.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<0>.MM_i_24_1 XI2.XI1.XI5.XI3<0>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<0>.MM_i_24_0 VDD! REG_DATA_9<0> XI2.XI1.XI5.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_9<0> XI2.XI1.XI5.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<0>.MM_i_24_1_48 XI2.XI1.XI5.XI3<0>.Y XI2.XI1.XI5.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<0>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<7>.MM_i_0 VSS! XI2.XI1.XI5.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<7>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<7>.MM_i_0_15 VSS! REG_DATA_9<7> XI2.XI1.XI5.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<7>.MM_i_0_15_63 XI2.XI1.XI5.XI3<7>.DUMMY1 REG_DATA_9<7>
+ XI2.XI1.XI5.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<7>.NEN
+ XI2.XI1.XI5.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<7>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<7>.MM_i_24 VDD! XI2.XI1.XI5.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<7>.MM_i_24_1 XI2.XI1.XI5.XI3<7>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<7>.MM_i_24_0 VDD! REG_DATA_9<7> XI2.XI1.XI5.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_9<7> XI2.XI1.XI5.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<7>.MM_i_24_1_48 XI2.XI1.XI5.XI3<7>.Y XI2.XI1.XI5.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<7>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<6>.MM_i_0 VSS! XI2.XI1.XI5.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<6>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<6>.MM_i_0_15 VSS! REG_DATA_9<6> XI2.XI1.XI5.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<6>.MM_i_0_15_63 XI2.XI1.XI5.XI3<6>.DUMMY1 REG_DATA_9<6>
+ XI2.XI1.XI5.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<6>.NEN
+ XI2.XI1.XI5.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<6>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<6>.MM_i_24 VDD! XI2.XI1.XI5.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<6>.MM_i_24_1 XI2.XI1.XI5.XI3<6>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<6>.MM_i_24_0 VDD! REG_DATA_9<6> XI2.XI1.XI5.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_9<6> XI2.XI1.XI5.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<6>.MM_i_24_1_48 XI2.XI1.XI5.XI3<6>.Y XI2.XI1.XI5.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<6>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<5>.MM_i_0 VSS! XI2.XI1.XI5.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<5>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<5>.MM_i_0_15 VSS! REG_DATA_9<5> XI2.XI1.XI5.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<5>.MM_i_0_15_63 XI2.XI1.XI5.XI3<5>.DUMMY1 REG_DATA_9<5>
+ XI2.XI1.XI5.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<5>.NEN
+ XI2.XI1.XI5.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<5>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<5>.MM_i_24 VDD! XI2.XI1.XI5.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<5>.MM_i_24_1 XI2.XI1.XI5.XI3<5>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<5>.MM_i_24_0 VDD! REG_DATA_9<5> XI2.XI1.XI5.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_9<5> XI2.XI1.XI5.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<5>.MM_i_24_1_48 XI2.XI1.XI5.XI3<5>.Y XI2.XI1.XI5.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<5>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<4>.MM_i_0 VSS! XI2.XI1.XI5.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<4>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<4>.MM_i_0_15 VSS! REG_DATA_9<4> XI2.XI1.XI5.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<4>.MM_i_0_15_63 XI2.XI1.XI5.XI3<4>.DUMMY1 REG_DATA_9<4>
+ XI2.XI1.XI5.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<4>.NEN
+ XI2.XI1.XI5.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<4>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<4>.MM_i_24 VDD! XI2.XI1.XI5.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<4>.MM_i_24_1 XI2.XI1.XI5.XI3<4>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<4>.MM_i_24_0 VDD! REG_DATA_9<4> XI2.XI1.XI5.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_9<4> XI2.XI1.XI5.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<4>.MM_i_24_1_48 XI2.XI1.XI5.XI3<4>.Y XI2.XI1.XI5.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<4>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<11>.MM_i_0 VSS! XI2.XI1.XI5.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<11>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<11>.MM_i_0_15 VSS! REG_DATA_9<11> XI2.XI1.XI5.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<11>.MM_i_0_15_63 XI2.XI1.XI5.XI3<11>.DUMMY1 REG_DATA_9<11>
+ XI2.XI1.XI5.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<11>.NEN
+ XI2.XI1.XI5.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<11>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<11>.MM_i_24 VDD! XI2.XI1.XI5.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<11>.MM_i_24_1 XI2.XI1.XI5.XI3<11>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<11>.MM_i_24_0 VDD! REG_DATA_9<11> XI2.XI1.XI5.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI5.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_9<11> XI2.XI1.XI5.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<11>.MM_i_24_1_48 XI2.XI1.XI5.XI3<11>.Y XI2.XI1.XI5.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<11>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<10>.MM_i_0 VSS! XI2.XI1.XI5.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<10>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<10>.MM_i_0_15 VSS! REG_DATA_9<10> XI2.XI1.XI5.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<10>.MM_i_0_15_63 XI2.XI1.XI5.XI3<10>.DUMMY1 REG_DATA_9<10>
+ XI2.XI1.XI5.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<10>.NEN
+ XI2.XI1.XI5.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<10>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<10>.MM_i_24 VDD! XI2.XI1.XI5.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<10>.MM_i_24_1 XI2.XI1.XI5.XI3<10>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<10>.MM_i_24_0 VDD! REG_DATA_9<10> XI2.XI1.XI5.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI5.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_9<10> XI2.XI1.XI5.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<10>.MM_i_24_1_48 XI2.XI1.XI5.XI3<10>.Y XI2.XI1.XI5.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<10>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<9>.MM_i_0 VSS! XI2.XI1.XI5.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<9>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<9>.MM_i_0_15 VSS! REG_DATA_9<9> XI2.XI1.XI5.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<9>.MM_i_0_15_63 XI2.XI1.XI5.XI3<9>.DUMMY1 REG_DATA_9<9>
+ XI2.XI1.XI5.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<9>.NEN
+ XI2.XI1.XI5.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<9>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<9>.MM_i_24 VDD! XI2.XI1.XI5.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<9>.MM_i_24_1 XI2.XI1.XI5.XI3<9>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<9>.MM_i_24_0 VDD! REG_DATA_9<9> XI2.XI1.XI5.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_9<9> XI2.XI1.XI5.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<9>.MM_i_24_1_48 XI2.XI1.XI5.XI3<9>.Y XI2.XI1.XI5.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<9>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<8>.MM_i_0 VSS! XI2.XI1.XI5.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<8>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<8>.MM_i_0_15 VSS! REG_DATA_9<8> XI2.XI1.XI5.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<8>.MM_i_0_15_63 XI2.XI1.XI5.XI3<8>.DUMMY1 REG_DATA_9<8>
+ XI2.XI1.XI5.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<8>.NEN
+ XI2.XI1.XI5.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<8>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<8>.MM_i_24 VDD! XI2.XI1.XI5.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<8>.MM_i_24_1 XI2.XI1.XI5.XI3<8>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<8>.MM_i_24_0 VDD! REG_DATA_9<8> XI2.XI1.XI5.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_9<8> XI2.XI1.XI5.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<8>.MM_i_24_1_48 XI2.XI1.XI5.XI3<8>.Y XI2.XI1.XI5.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<8>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<15>.MM_i_0 VSS! XI2.XI1.XI5.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<15>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<15>.MM_i_0_15 VSS! REG_DATA_9<15> XI2.XI1.XI5.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<15>.MM_i_0_15_63 XI2.XI1.XI5.XI3<15>.DUMMY1 REG_DATA_9<15>
+ XI2.XI1.XI5.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<15>.NEN
+ XI2.XI1.XI5.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<15>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<15>.MM_i_24 VDD! XI2.XI1.XI5.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<15>.MM_i_24_1 XI2.XI1.XI5.XI3<15>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<15>.MM_i_24_0 VDD! REG_DATA_9<15> XI2.XI1.XI5.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI5.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_9<15> XI2.XI1.XI5.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<15>.MM_i_24_1_48 XI2.XI1.XI5.XI3<15>.Y XI2.XI1.XI5.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<15>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<14>.MM_i_0 VSS! XI2.XI1.XI5.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<14>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<14>.MM_i_0_15 VSS! REG_DATA_9<14> XI2.XI1.XI5.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<14>.MM_i_0_15_63 XI2.XI1.XI5.XI3<14>.DUMMY1 REG_DATA_9<14>
+ XI2.XI1.XI5.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<14>.NEN
+ XI2.XI1.XI5.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<14>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<14>.MM_i_24 VDD! XI2.XI1.XI5.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<14>.MM_i_24_1 XI2.XI1.XI5.XI3<14>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<14>.MM_i_24_0 VDD! REG_DATA_9<14> XI2.XI1.XI5.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI5.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_9<14> XI2.XI1.XI5.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<14>.MM_i_24_1_48 XI2.XI1.XI5.XI3<14>.Y XI2.XI1.XI5.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<14>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<13>.MM_i_0 VSS! XI2.XI1.XI5.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<13>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<13>.MM_i_0_15 VSS! REG_DATA_9<13> XI2.XI1.XI5.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<13>.MM_i_0_15_63 XI2.XI1.XI5.XI3<13>.DUMMY1 REG_DATA_9<13>
+ XI2.XI1.XI5.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<13>.NEN
+ XI2.XI1.XI5.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<13>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<13>.MM_i_24 VDD! XI2.XI1.XI5.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<13>.MM_i_24_1 XI2.XI1.XI5.XI3<13>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<13>.MM_i_24_0 VDD! REG_DATA_9<13> XI2.XI1.XI5.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI5.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_9<13> XI2.XI1.XI5.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<13>.MM_i_24_1_48 XI2.XI1.XI5.XI3<13>.Y XI2.XI1.XI5.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<13>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI5.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI5.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI5.XI3<12>.MM_i_0 VSS! XI2.XI1.XI5.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI5.XI3<12>.MM_i_0_14 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<12>.MM_i_0_15 VSS! REG_DATA_9<12> XI2.XI1.XI5.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<12>.MM_i_0_15_63 XI2.XI1.XI5.XI3<12>.DUMMY1 REG_DATA_9<12>
+ XI2.XI1.XI5.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI5.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI5.XI3<12>.NEN
+ XI2.XI1.XI5.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI5.XI3<12>.MM_i_17 VSS! XI2.NET1<3> XI2.XI1.XI5.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI5.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI5.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<12>.MM_i_24 VDD! XI2.XI1.XI5.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI5.XI3<12>.MM_i_24_1 XI2.XI1.XI5.XI3<12>.DUMMY0 XI2.NET1<3>
+ XI2.XI1.XI5.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI5.XI3<12>.MM_i_24_0 VDD! REG_DATA_9<12> XI2.XI1.XI5.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI5.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_9<12> XI2.XI1.XI5.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI5.XI3<12>.MM_i_24_1_48 XI2.XI1.XI5.XI3<12>.Y XI2.XI1.XI5.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI5.XI3<12>.MM_i_42 VDD! XI2.NET1<3> XI2.XI1.XI5.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<3>.MM_i_0 VSS! XI2.XI1.XI10.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<3>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<3>.MM_i_0_15 VSS! REG_DATA_8<3> XI2.XI1.XI10.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<3>.MM_i_0_15_63 XI2.XI1.XI10.XI3<3>.DUMMY1 REG_DATA_8<3>
+ XI2.XI1.XI10.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<3>.NEN
+ XI2.XI1.XI10.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<3>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<3>.MM_i_24 VDD! XI2.XI1.XI10.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<3>.MM_i_24_1 XI2.XI1.XI10.XI3<3>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<3>.MM_i_24_0 VDD! REG_DATA_8<3> XI2.XI1.XI10.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_8<3> XI2.XI1.XI10.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<3>.MM_i_24_1_48 XI2.XI1.XI10.XI3<3>.Y XI2.XI1.XI10.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<3>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<2>.MM_i_0 VSS! XI2.XI1.XI10.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<2>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<2>.MM_i_0_15 VSS! REG_DATA_8<2> XI2.XI1.XI10.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<2>.MM_i_0_15_63 XI2.XI1.XI10.XI3<2>.DUMMY1 REG_DATA_8<2>
+ XI2.XI1.XI10.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<2>.NEN
+ XI2.XI1.XI10.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<2>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<2>.MM_i_24 VDD! XI2.XI1.XI10.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<2>.MM_i_24_1 XI2.XI1.XI10.XI3<2>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<2>.MM_i_24_0 VDD! REG_DATA_8<2> XI2.XI1.XI10.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_8<2> XI2.XI1.XI10.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<2>.MM_i_24_1_48 XI2.XI1.XI10.XI3<2>.Y XI2.XI1.XI10.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<2>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<1>.MM_i_0 VSS! XI2.XI1.XI10.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<1>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<1>.MM_i_0_15 VSS! REG_DATA_8<1> XI2.XI1.XI10.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<1>.MM_i_0_15_63 XI2.XI1.XI10.XI3<1>.DUMMY1 REG_DATA_8<1>
+ XI2.XI1.XI10.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<1>.NEN
+ XI2.XI1.XI10.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<1>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<1>.MM_i_24 VDD! XI2.XI1.XI10.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<1>.MM_i_24_1 XI2.XI1.XI10.XI3<1>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<1>.MM_i_24_0 VDD! REG_DATA_8<1> XI2.XI1.XI10.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_8<1> XI2.XI1.XI10.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<1>.MM_i_24_1_48 XI2.XI1.XI10.XI3<1>.Y XI2.XI1.XI10.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<1>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<0>.MM_i_0 VSS! XI2.XI1.XI10.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<0>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<0>.MM_i_0_15 VSS! REG_DATA_8<0> XI2.XI1.XI10.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<0>.MM_i_0_15_63 XI2.XI1.XI10.XI3<0>.DUMMY1 REG_DATA_8<0>
+ XI2.XI1.XI10.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<0>.NEN
+ XI2.XI1.XI10.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<0>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<0>.MM_i_24 VDD! XI2.XI1.XI10.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<0>.MM_i_24_1 XI2.XI1.XI10.XI3<0>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<0>.MM_i_24_0 VDD! REG_DATA_8<0> XI2.XI1.XI10.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_8<0> XI2.XI1.XI10.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<0>.MM_i_24_1_48 XI2.XI1.XI10.XI3<0>.Y XI2.XI1.XI10.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<0>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<7>.MM_i_0 VSS! XI2.XI1.XI10.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<7>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<7>.MM_i_0_15 VSS! REG_DATA_8<7> XI2.XI1.XI10.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<7>.MM_i_0_15_63 XI2.XI1.XI10.XI3<7>.DUMMY1 REG_DATA_8<7>
+ XI2.XI1.XI10.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<7>.NEN
+ XI2.XI1.XI10.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<7>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<7>.MM_i_24 VDD! XI2.XI1.XI10.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<7>.MM_i_24_1 XI2.XI1.XI10.XI3<7>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<7>.MM_i_24_0 VDD! REG_DATA_8<7> XI2.XI1.XI10.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_8<7> XI2.XI1.XI10.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<7>.MM_i_24_1_48 XI2.XI1.XI10.XI3<7>.Y XI2.XI1.XI10.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<7>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<6>.MM_i_0 VSS! XI2.XI1.XI10.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<6>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<6>.MM_i_0_15 VSS! REG_DATA_8<6> XI2.XI1.XI10.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<6>.MM_i_0_15_63 XI2.XI1.XI10.XI3<6>.DUMMY1 REG_DATA_8<6>
+ XI2.XI1.XI10.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<6>.NEN
+ XI2.XI1.XI10.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<6>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<6>.MM_i_24 VDD! XI2.XI1.XI10.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<6>.MM_i_24_1 XI2.XI1.XI10.XI3<6>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<6>.MM_i_24_0 VDD! REG_DATA_8<6> XI2.XI1.XI10.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_8<6> XI2.XI1.XI10.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<6>.MM_i_24_1_48 XI2.XI1.XI10.XI3<6>.Y XI2.XI1.XI10.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<6>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<5>.MM_i_0 VSS! XI2.XI1.XI10.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<5>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<5>.MM_i_0_15 VSS! REG_DATA_8<5> XI2.XI1.XI10.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<5>.MM_i_0_15_63 XI2.XI1.XI10.XI3<5>.DUMMY1 REG_DATA_8<5>
+ XI2.XI1.XI10.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<5>.NEN
+ XI2.XI1.XI10.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<5>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<5>.MM_i_24 VDD! XI2.XI1.XI10.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<5>.MM_i_24_1 XI2.XI1.XI10.XI3<5>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<5>.MM_i_24_0 VDD! REG_DATA_8<5> XI2.XI1.XI10.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_8<5> XI2.XI1.XI10.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<5>.MM_i_24_1_48 XI2.XI1.XI10.XI3<5>.Y XI2.XI1.XI10.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<5>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<4>.MM_i_0 VSS! XI2.XI1.XI10.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<4>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<4>.MM_i_0_15 VSS! REG_DATA_8<4> XI2.XI1.XI10.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<4>.MM_i_0_15_63 XI2.XI1.XI10.XI3<4>.DUMMY1 REG_DATA_8<4>
+ XI2.XI1.XI10.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<4>.NEN
+ XI2.XI1.XI10.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<4>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<4>.MM_i_24 VDD! XI2.XI1.XI10.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<4>.MM_i_24_1 XI2.XI1.XI10.XI3<4>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<4>.MM_i_24_0 VDD! REG_DATA_8<4> XI2.XI1.XI10.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_8<4> XI2.XI1.XI10.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<4>.MM_i_24_1_48 XI2.XI1.XI10.XI3<4>.Y XI2.XI1.XI10.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<4>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<11>.MM_i_0 VSS! XI2.XI1.XI10.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<11>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<11>.MM_i_0_15 VSS! REG_DATA_8<11> XI2.XI1.XI10.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<11>.MM_i_0_15_63 XI2.XI1.XI10.XI3<11>.DUMMY1 REG_DATA_8<11>
+ XI2.XI1.XI10.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<11>.NEN
+ XI2.XI1.XI10.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<11>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<11>.MM_i_24 VDD! XI2.XI1.XI10.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<11>.MM_i_24_1 XI2.XI1.XI10.XI3<11>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<11>.MM_i_24_0 VDD! REG_DATA_8<11> XI2.XI1.XI10.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_8<11> XI2.XI1.XI10.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<11>.MM_i_24_1_48 XI2.XI1.XI10.XI3<11>.Y
+ XI2.XI1.XI10.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI10.XI3<11>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<10>.MM_i_0 VSS! XI2.XI1.XI10.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<10>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<10>.MM_i_0_15 VSS! REG_DATA_8<10> XI2.XI1.XI10.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<10>.MM_i_0_15_63 XI2.XI1.XI10.XI3<10>.DUMMY1 REG_DATA_8<10>
+ XI2.XI1.XI10.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<10>.NEN
+ XI2.XI1.XI10.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<10>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<10>.MM_i_24 VDD! XI2.XI1.XI10.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<10>.MM_i_24_1 XI2.XI1.XI10.XI3<10>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<10>.MM_i_24_0 VDD! REG_DATA_8<10> XI2.XI1.XI10.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_8<10> XI2.XI1.XI10.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<10>.MM_i_24_1_48 XI2.XI1.XI10.XI3<10>.Y
+ XI2.XI1.XI10.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI10.XI3<10>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<9>.MM_i_0 VSS! XI2.XI1.XI10.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<9>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<9>.MM_i_0_15 VSS! REG_DATA_8<9> XI2.XI1.XI10.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<9>.MM_i_0_15_63 XI2.XI1.XI10.XI3<9>.DUMMY1 REG_DATA_8<9>
+ XI2.XI1.XI10.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<9>.NEN
+ XI2.XI1.XI10.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<9>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<9>.MM_i_24 VDD! XI2.XI1.XI10.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<9>.MM_i_24_1 XI2.XI1.XI10.XI3<9>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<9>.MM_i_24_0 VDD! REG_DATA_8<9> XI2.XI1.XI10.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_8<9> XI2.XI1.XI10.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<9>.MM_i_24_1_48 XI2.XI1.XI10.XI3<9>.Y XI2.XI1.XI10.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<9>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<8>.MM_i_0 VSS! XI2.XI1.XI10.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<8>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<8>.MM_i_0_15 VSS! REG_DATA_8<8> XI2.XI1.XI10.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<8>.MM_i_0_15_63 XI2.XI1.XI10.XI3<8>.DUMMY1 REG_DATA_8<8>
+ XI2.XI1.XI10.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<8>.NEN
+ XI2.XI1.XI10.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<8>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<8>.MM_i_24 VDD! XI2.XI1.XI10.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<8>.MM_i_24_1 XI2.XI1.XI10.XI3<8>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<8>.MM_i_24_0 VDD! REG_DATA_8<8> XI2.XI1.XI10.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_8<8> XI2.XI1.XI10.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI10.XI3<8>.MM_i_24_1_48 XI2.XI1.XI10.XI3<8>.Y XI2.XI1.XI10.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI10.XI3<8>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<15>.MM_i_0 VSS! XI2.XI1.XI10.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<15>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<15>.MM_i_0_15 VSS! REG_DATA_8<15> XI2.XI1.XI10.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<15>.MM_i_0_15_63 XI2.XI1.XI10.XI3<15>.DUMMY1 REG_DATA_8<15>
+ XI2.XI1.XI10.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<15>.NEN
+ XI2.XI1.XI10.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<15>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<15>.MM_i_24 VDD! XI2.XI1.XI10.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<15>.MM_i_24_1 XI2.XI1.XI10.XI3<15>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<15>.MM_i_24_0 VDD! REG_DATA_8<15> XI2.XI1.XI10.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_8<15> XI2.XI1.XI10.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<15>.MM_i_24_1_48 XI2.XI1.XI10.XI3<15>.Y
+ XI2.XI1.XI10.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI10.XI3<15>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<14>.MM_i_0 VSS! XI2.XI1.XI10.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<14>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<14>.MM_i_0_15 VSS! REG_DATA_8<14> XI2.XI1.XI10.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<14>.MM_i_0_15_63 XI2.XI1.XI10.XI3<14>.DUMMY1 REG_DATA_8<14>
+ XI2.XI1.XI10.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<14>.NEN
+ XI2.XI1.XI10.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<14>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<14>.MM_i_24 VDD! XI2.XI1.XI10.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<14>.MM_i_24_1 XI2.XI1.XI10.XI3<14>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<14>.MM_i_24_0 VDD! REG_DATA_8<14> XI2.XI1.XI10.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_8<14> XI2.XI1.XI10.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<14>.MM_i_24_1_48 XI2.XI1.XI10.XI3<14>.Y
+ XI2.XI1.XI10.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI10.XI3<14>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<13>.MM_i_0 VSS! XI2.XI1.XI10.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<13>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<13>.MM_i_0_15 VSS! REG_DATA_8<13> XI2.XI1.XI10.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<13>.MM_i_0_15_63 XI2.XI1.XI10.XI3<13>.DUMMY1 REG_DATA_8<13>
+ XI2.XI1.XI10.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<13>.NEN
+ XI2.XI1.XI10.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<13>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<13>.MM_i_24 VDD! XI2.XI1.XI10.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<13>.MM_i_24_1 XI2.XI1.XI10.XI3<13>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<13>.MM_i_24_0 VDD! REG_DATA_8<13> XI2.XI1.XI10.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_8<13> XI2.XI1.XI10.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<13>.MM_i_24_1_48 XI2.XI1.XI10.XI3<13>.Y
+ XI2.XI1.XI10.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI10.XI3<13>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI10.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI10.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI10.XI3<12>.MM_i_0 VSS! XI2.XI1.XI10.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI10.XI3<12>.MM_i_0_14 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<12>.MM_i_0_15 VSS! REG_DATA_8<12> XI2.XI1.XI10.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<12>.MM_i_0_15_63 XI2.XI1.XI10.XI3<12>.DUMMY1 REG_DATA_8<12>
+ XI2.XI1.XI10.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI10.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI10.XI3<12>.NEN
+ XI2.XI1.XI10.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI10.XI3<12>.MM_i_17 VSS! XI2.NET1<4> XI2.XI1.XI10.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI10.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI10.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<12>.MM_i_24 VDD! XI2.XI1.XI10.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI10.XI3<12>.MM_i_24_1 XI2.XI1.XI10.XI3<12>.DUMMY0 XI2.NET1<4>
+ XI2.XI1.XI10.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI10.XI3<12>.MM_i_24_0 VDD! REG_DATA_8<12> XI2.XI1.XI10.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_8<12> XI2.XI1.XI10.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI10.XI3<12>.MM_i_24_1_48 XI2.XI1.XI10.XI3<12>.Y
+ XI2.XI1.XI10.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI10.XI3<12>.MM_i_42 VDD! XI2.NET1<4> XI2.XI1.XI10.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<3>.MM_i_0 VSS! XI2.XI1.XI9.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<3>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<3>.MM_i_0_15 VSS! REG_DATA_7<3> XI2.XI1.XI9.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<3>.MM_i_0_15_63 XI2.XI1.XI9.XI3<3>.DUMMY1 REG_DATA_7<3>
+ XI2.XI1.XI9.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<3>.NEN
+ XI2.XI1.XI9.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<3>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<3>.MM_i_24 VDD! XI2.XI1.XI9.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<3>.MM_i_24_1 XI2.XI1.XI9.XI3<3>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<3>.MM_i_24_0 VDD! REG_DATA_7<3> XI2.XI1.XI9.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_7<3> XI2.XI1.XI9.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<3>.MM_i_24_1_48 XI2.XI1.XI9.XI3<3>.Y XI2.XI1.XI9.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<3>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<2>.MM_i_0 VSS! XI2.XI1.XI9.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<2>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<2>.MM_i_0_15 VSS! REG_DATA_7<2> XI2.XI1.XI9.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<2>.MM_i_0_15_63 XI2.XI1.XI9.XI3<2>.DUMMY1 REG_DATA_7<2>
+ XI2.XI1.XI9.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<2>.NEN
+ XI2.XI1.XI9.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<2>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<2>.MM_i_24 VDD! XI2.XI1.XI9.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<2>.MM_i_24_1 XI2.XI1.XI9.XI3<2>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<2>.MM_i_24_0 VDD! REG_DATA_7<2> XI2.XI1.XI9.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_7<2> XI2.XI1.XI9.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<2>.MM_i_24_1_48 XI2.XI1.XI9.XI3<2>.Y XI2.XI1.XI9.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<2>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<1>.MM_i_0 VSS! XI2.XI1.XI9.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<1>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<1>.MM_i_0_15 VSS! REG_DATA_7<1> XI2.XI1.XI9.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<1>.MM_i_0_15_63 XI2.XI1.XI9.XI3<1>.DUMMY1 REG_DATA_7<1>
+ XI2.XI1.XI9.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<1>.NEN
+ XI2.XI1.XI9.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<1>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<1>.MM_i_24 VDD! XI2.XI1.XI9.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<1>.MM_i_24_1 XI2.XI1.XI9.XI3<1>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<1>.MM_i_24_0 VDD! REG_DATA_7<1> XI2.XI1.XI9.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_7<1> XI2.XI1.XI9.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<1>.MM_i_24_1_48 XI2.XI1.XI9.XI3<1>.Y XI2.XI1.XI9.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<1>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<0>.MM_i_0 VSS! XI2.XI1.XI9.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<0>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<0>.MM_i_0_15 VSS! REG_DATA_7<0> XI2.XI1.XI9.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<0>.MM_i_0_15_63 XI2.XI1.XI9.XI3<0>.DUMMY1 REG_DATA_7<0>
+ XI2.XI1.XI9.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<0>.NEN
+ XI2.XI1.XI9.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<0>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<0>.MM_i_24 VDD! XI2.XI1.XI9.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<0>.MM_i_24_1 XI2.XI1.XI9.XI3<0>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<0>.MM_i_24_0 VDD! REG_DATA_7<0> XI2.XI1.XI9.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_7<0> XI2.XI1.XI9.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<0>.MM_i_24_1_48 XI2.XI1.XI9.XI3<0>.Y XI2.XI1.XI9.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<0>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<7>.MM_i_0 VSS! XI2.XI1.XI9.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<7>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<7>.MM_i_0_15 VSS! REG_DATA_7<7> XI2.XI1.XI9.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<7>.MM_i_0_15_63 XI2.XI1.XI9.XI3<7>.DUMMY1 REG_DATA_7<7>
+ XI2.XI1.XI9.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<7>.NEN
+ XI2.XI1.XI9.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<7>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<7>.MM_i_24 VDD! XI2.XI1.XI9.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<7>.MM_i_24_1 XI2.XI1.XI9.XI3<7>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<7>.MM_i_24_0 VDD! REG_DATA_7<7> XI2.XI1.XI9.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_7<7> XI2.XI1.XI9.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<7>.MM_i_24_1_48 XI2.XI1.XI9.XI3<7>.Y XI2.XI1.XI9.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<7>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<6>.MM_i_0 VSS! XI2.XI1.XI9.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<6>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<6>.MM_i_0_15 VSS! REG_DATA_7<6> XI2.XI1.XI9.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<6>.MM_i_0_15_63 XI2.XI1.XI9.XI3<6>.DUMMY1 REG_DATA_7<6>
+ XI2.XI1.XI9.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<6>.NEN
+ XI2.XI1.XI9.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<6>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<6>.MM_i_24 VDD! XI2.XI1.XI9.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<6>.MM_i_24_1 XI2.XI1.XI9.XI3<6>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<6>.MM_i_24_0 VDD! REG_DATA_7<6> XI2.XI1.XI9.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_7<6> XI2.XI1.XI9.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<6>.MM_i_24_1_48 XI2.XI1.XI9.XI3<6>.Y XI2.XI1.XI9.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<6>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<5>.MM_i_0 VSS! XI2.XI1.XI9.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<5>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<5>.MM_i_0_15 VSS! REG_DATA_7<5> XI2.XI1.XI9.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<5>.MM_i_0_15_63 XI2.XI1.XI9.XI3<5>.DUMMY1 REG_DATA_7<5>
+ XI2.XI1.XI9.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<5>.NEN
+ XI2.XI1.XI9.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<5>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<5>.MM_i_24 VDD! XI2.XI1.XI9.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<5>.MM_i_24_1 XI2.XI1.XI9.XI3<5>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<5>.MM_i_24_0 VDD! REG_DATA_7<5> XI2.XI1.XI9.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_7<5> XI2.XI1.XI9.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<5>.MM_i_24_1_48 XI2.XI1.XI9.XI3<5>.Y XI2.XI1.XI9.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<5>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<4>.MM_i_0 VSS! XI2.XI1.XI9.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<4>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<4>.MM_i_0_15 VSS! REG_DATA_7<4> XI2.XI1.XI9.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<4>.MM_i_0_15_63 XI2.XI1.XI9.XI3<4>.DUMMY1 REG_DATA_7<4>
+ XI2.XI1.XI9.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<4>.NEN
+ XI2.XI1.XI9.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<4>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<4>.MM_i_24 VDD! XI2.XI1.XI9.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<4>.MM_i_24_1 XI2.XI1.XI9.XI3<4>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<4>.MM_i_24_0 VDD! REG_DATA_7<4> XI2.XI1.XI9.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_7<4> XI2.XI1.XI9.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<4>.MM_i_24_1_48 XI2.XI1.XI9.XI3<4>.Y XI2.XI1.XI9.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<4>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<11>.MM_i_0 VSS! XI2.XI1.XI9.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<11>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<11>.MM_i_0_15 VSS! REG_DATA_7<11> XI2.XI1.XI9.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<11>.MM_i_0_15_63 XI2.XI1.XI9.XI3<11>.DUMMY1 REG_DATA_7<11>
+ XI2.XI1.XI9.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<11>.NEN
+ XI2.XI1.XI9.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<11>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<11>.MM_i_24 VDD! XI2.XI1.XI9.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<11>.MM_i_24_1 XI2.XI1.XI9.XI3<11>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<11>.MM_i_24_0 VDD! REG_DATA_7<11> XI2.XI1.XI9.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI9.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_7<11> XI2.XI1.XI9.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<11>.MM_i_24_1_48 XI2.XI1.XI9.XI3<11>.Y XI2.XI1.XI9.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<11>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<10>.MM_i_0 VSS! XI2.XI1.XI9.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<10>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<10>.MM_i_0_15 VSS! REG_DATA_7<10> XI2.XI1.XI9.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<10>.MM_i_0_15_63 XI2.XI1.XI9.XI3<10>.DUMMY1 REG_DATA_7<10>
+ XI2.XI1.XI9.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<10>.NEN
+ XI2.XI1.XI9.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<10>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<10>.MM_i_24 VDD! XI2.XI1.XI9.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<10>.MM_i_24_1 XI2.XI1.XI9.XI3<10>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<10>.MM_i_24_0 VDD! REG_DATA_7<10> XI2.XI1.XI9.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI9.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_7<10> XI2.XI1.XI9.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<10>.MM_i_24_1_48 XI2.XI1.XI9.XI3<10>.Y XI2.XI1.XI9.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<10>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<9>.MM_i_0 VSS! XI2.XI1.XI9.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<9>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<9>.MM_i_0_15 VSS! REG_DATA_7<9> XI2.XI1.XI9.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<9>.MM_i_0_15_63 XI2.XI1.XI9.XI3<9>.DUMMY1 REG_DATA_7<9>
+ XI2.XI1.XI9.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<9>.NEN
+ XI2.XI1.XI9.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<9>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<9>.MM_i_24 VDD! XI2.XI1.XI9.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<9>.MM_i_24_1 XI2.XI1.XI9.XI3<9>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<9>.MM_i_24_0 VDD! REG_DATA_7<9> XI2.XI1.XI9.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_7<9> XI2.XI1.XI9.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<9>.MM_i_24_1_48 XI2.XI1.XI9.XI3<9>.Y XI2.XI1.XI9.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<9>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<8>.MM_i_0 VSS! XI2.XI1.XI9.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<8>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<8>.MM_i_0_15 VSS! REG_DATA_7<8> XI2.XI1.XI9.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<8>.MM_i_0_15_63 XI2.XI1.XI9.XI3<8>.DUMMY1 REG_DATA_7<8>
+ XI2.XI1.XI9.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<8>.NEN
+ XI2.XI1.XI9.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<8>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<8>.MM_i_24 VDD! XI2.XI1.XI9.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<8>.MM_i_24_1 XI2.XI1.XI9.XI3<8>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<8>.MM_i_24_0 VDD! REG_DATA_7<8> XI2.XI1.XI9.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_7<8> XI2.XI1.XI9.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<8>.MM_i_24_1_48 XI2.XI1.XI9.XI3<8>.Y XI2.XI1.XI9.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<8>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<15>.MM_i_0 VSS! XI2.XI1.XI9.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<15>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<15>.MM_i_0_15 VSS! REG_DATA_7<15> XI2.XI1.XI9.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<15>.MM_i_0_15_63 XI2.XI1.XI9.XI3<15>.DUMMY1 REG_DATA_7<15>
+ XI2.XI1.XI9.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<15>.NEN
+ XI2.XI1.XI9.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<15>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<15>.MM_i_24 VDD! XI2.XI1.XI9.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<15>.MM_i_24_1 XI2.XI1.XI9.XI3<15>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<15>.MM_i_24_0 VDD! REG_DATA_7<15> XI2.XI1.XI9.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI9.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_7<15> XI2.XI1.XI9.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<15>.MM_i_24_1_48 XI2.XI1.XI9.XI3<15>.Y XI2.XI1.XI9.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<15>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<14>.MM_i_0 VSS! XI2.XI1.XI9.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<14>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<14>.MM_i_0_15 VSS! REG_DATA_7<14> XI2.XI1.XI9.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<14>.MM_i_0_15_63 XI2.XI1.XI9.XI3<14>.DUMMY1 REG_DATA_7<14>
+ XI2.XI1.XI9.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<14>.NEN
+ XI2.XI1.XI9.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<14>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<14>.MM_i_24 VDD! XI2.XI1.XI9.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<14>.MM_i_24_1 XI2.XI1.XI9.XI3<14>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<14>.MM_i_24_0 VDD! REG_DATA_7<14> XI2.XI1.XI9.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI9.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_7<14> XI2.XI1.XI9.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<14>.MM_i_24_1_48 XI2.XI1.XI9.XI3<14>.Y XI2.XI1.XI9.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<14>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<13>.MM_i_0 VSS! XI2.XI1.XI9.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<13>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<13>.MM_i_0_15 VSS! REG_DATA_7<13> XI2.XI1.XI9.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<13>.MM_i_0_15_63 XI2.XI1.XI9.XI3<13>.DUMMY1 REG_DATA_7<13>
+ XI2.XI1.XI9.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<13>.NEN
+ XI2.XI1.XI9.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<13>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<13>.MM_i_24 VDD! XI2.XI1.XI9.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<13>.MM_i_24_1 XI2.XI1.XI9.XI3<13>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<13>.MM_i_24_0 VDD! REG_DATA_7<13> XI2.XI1.XI9.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI9.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_7<13> XI2.XI1.XI9.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<13>.MM_i_24_1_48 XI2.XI1.XI9.XI3<13>.Y XI2.XI1.XI9.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<13>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI9.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI9.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI9.XI3<12>.MM_i_0 VSS! XI2.XI1.XI9.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI9.XI3<12>.MM_i_0_14 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<12>.MM_i_0_15 VSS! REG_DATA_7<12> XI2.XI1.XI9.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<12>.MM_i_0_15_63 XI2.XI1.XI9.XI3<12>.DUMMY1 REG_DATA_7<12>
+ XI2.XI1.XI9.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI9.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI9.XI3<12>.NEN
+ XI2.XI1.XI9.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI9.XI3<12>.MM_i_17 VSS! XI2.NET1<5> XI2.XI1.XI9.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI9.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI9.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<12>.MM_i_24 VDD! XI2.XI1.XI9.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI9.XI3<12>.MM_i_24_1 XI2.XI1.XI9.XI3<12>.DUMMY0 XI2.NET1<5>
+ XI2.XI1.XI9.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI9.XI3<12>.MM_i_24_0 VDD! REG_DATA_7<12> XI2.XI1.XI9.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI9.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_7<12> XI2.XI1.XI9.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI9.XI3<12>.MM_i_24_1_48 XI2.XI1.XI9.XI3<12>.Y XI2.XI1.XI9.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI9.XI3<12>.MM_i_42 VDD! XI2.NET1<5> XI2.XI1.XI9.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<3>.MM_i_0 VSS! XI2.XI1.XI7.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<3>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<3>.MM_i_0_15 VSS! REG_DATA_6<3> XI2.XI1.XI7.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<3>.MM_i_0_15_63 XI2.XI1.XI7.XI3<3>.DUMMY1 REG_DATA_6<3>
+ XI2.XI1.XI7.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<3>.NEN
+ XI2.XI1.XI7.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<3>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<3>.MM_i_24 VDD! XI2.XI1.XI7.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<3>.MM_i_24_1 XI2.XI1.XI7.XI3<3>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<3>.MM_i_24_0 VDD! REG_DATA_6<3> XI2.XI1.XI7.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_6<3> XI2.XI1.XI7.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<3>.MM_i_24_1_48 XI2.XI1.XI7.XI3<3>.Y XI2.XI1.XI7.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<3>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<2>.MM_i_0 VSS! XI2.XI1.XI7.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<2>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<2>.MM_i_0_15 VSS! REG_DATA_6<2> XI2.XI1.XI7.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<2>.MM_i_0_15_63 XI2.XI1.XI7.XI3<2>.DUMMY1 REG_DATA_6<2>
+ XI2.XI1.XI7.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<2>.NEN
+ XI2.XI1.XI7.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<2>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<2>.MM_i_24 VDD! XI2.XI1.XI7.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<2>.MM_i_24_1 XI2.XI1.XI7.XI3<2>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<2>.MM_i_24_0 VDD! REG_DATA_6<2> XI2.XI1.XI7.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_6<2> XI2.XI1.XI7.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<2>.MM_i_24_1_48 XI2.XI1.XI7.XI3<2>.Y XI2.XI1.XI7.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<2>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<1>.MM_i_0 VSS! XI2.XI1.XI7.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<1>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<1>.MM_i_0_15 VSS! REG_DATA_6<1> XI2.XI1.XI7.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<1>.MM_i_0_15_63 XI2.XI1.XI7.XI3<1>.DUMMY1 REG_DATA_6<1>
+ XI2.XI1.XI7.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<1>.NEN
+ XI2.XI1.XI7.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<1>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<1>.MM_i_24 VDD! XI2.XI1.XI7.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<1>.MM_i_24_1 XI2.XI1.XI7.XI3<1>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<1>.MM_i_24_0 VDD! REG_DATA_6<1> XI2.XI1.XI7.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_6<1> XI2.XI1.XI7.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<1>.MM_i_24_1_48 XI2.XI1.XI7.XI3<1>.Y XI2.XI1.XI7.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<1>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<0>.MM_i_0 VSS! XI2.XI1.XI7.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<0>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<0>.MM_i_0_15 VSS! REG_DATA_6<0> XI2.XI1.XI7.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<0>.MM_i_0_15_63 XI2.XI1.XI7.XI3<0>.DUMMY1 REG_DATA_6<0>
+ XI2.XI1.XI7.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<0>.NEN
+ XI2.XI1.XI7.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<0>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<0>.MM_i_24 VDD! XI2.XI1.XI7.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<0>.MM_i_24_1 XI2.XI1.XI7.XI3<0>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<0>.MM_i_24_0 VDD! REG_DATA_6<0> XI2.XI1.XI7.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_6<0> XI2.XI1.XI7.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<0>.MM_i_24_1_48 XI2.XI1.XI7.XI3<0>.Y XI2.XI1.XI7.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<0>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<7>.MM_i_0 VSS! XI2.XI1.XI7.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<7>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<7>.MM_i_0_15 VSS! REG_DATA_6<7> XI2.XI1.XI7.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<7>.MM_i_0_15_63 XI2.XI1.XI7.XI3<7>.DUMMY1 REG_DATA_6<7>
+ XI2.XI1.XI7.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<7>.NEN
+ XI2.XI1.XI7.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<7>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<7>.MM_i_24 VDD! XI2.XI1.XI7.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<7>.MM_i_24_1 XI2.XI1.XI7.XI3<7>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<7>.MM_i_24_0 VDD! REG_DATA_6<7> XI2.XI1.XI7.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_6<7> XI2.XI1.XI7.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<7>.MM_i_24_1_48 XI2.XI1.XI7.XI3<7>.Y XI2.XI1.XI7.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<7>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<6>.MM_i_0 VSS! XI2.XI1.XI7.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<6>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<6>.MM_i_0_15 VSS! REG_DATA_6<6> XI2.XI1.XI7.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<6>.MM_i_0_15_63 XI2.XI1.XI7.XI3<6>.DUMMY1 REG_DATA_6<6>
+ XI2.XI1.XI7.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<6>.NEN
+ XI2.XI1.XI7.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<6>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<6>.MM_i_24 VDD! XI2.XI1.XI7.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<6>.MM_i_24_1 XI2.XI1.XI7.XI3<6>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<6>.MM_i_24_0 VDD! REG_DATA_6<6> XI2.XI1.XI7.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_6<6> XI2.XI1.XI7.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<6>.MM_i_24_1_48 XI2.XI1.XI7.XI3<6>.Y XI2.XI1.XI7.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<6>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<5>.MM_i_0 VSS! XI2.XI1.XI7.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<5>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<5>.MM_i_0_15 VSS! REG_DATA_6<5> XI2.XI1.XI7.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<5>.MM_i_0_15_63 XI2.XI1.XI7.XI3<5>.DUMMY1 REG_DATA_6<5>
+ XI2.XI1.XI7.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<5>.NEN
+ XI2.XI1.XI7.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<5>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<5>.MM_i_24 VDD! XI2.XI1.XI7.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<5>.MM_i_24_1 XI2.XI1.XI7.XI3<5>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<5>.MM_i_24_0 VDD! REG_DATA_6<5> XI2.XI1.XI7.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_6<5> XI2.XI1.XI7.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<5>.MM_i_24_1_48 XI2.XI1.XI7.XI3<5>.Y XI2.XI1.XI7.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<5>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<4>.MM_i_0 VSS! XI2.XI1.XI7.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<4>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<4>.MM_i_0_15 VSS! REG_DATA_6<4> XI2.XI1.XI7.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<4>.MM_i_0_15_63 XI2.XI1.XI7.XI3<4>.DUMMY1 REG_DATA_6<4>
+ XI2.XI1.XI7.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<4>.NEN
+ XI2.XI1.XI7.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<4>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<4>.MM_i_24 VDD! XI2.XI1.XI7.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<4>.MM_i_24_1 XI2.XI1.XI7.XI3<4>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<4>.MM_i_24_0 VDD! REG_DATA_6<4> XI2.XI1.XI7.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_6<4> XI2.XI1.XI7.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<4>.MM_i_24_1_48 XI2.XI1.XI7.XI3<4>.Y XI2.XI1.XI7.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<4>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<11>.MM_i_0 VSS! XI2.XI1.XI7.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<11>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<11>.MM_i_0_15 VSS! REG_DATA_6<11> XI2.XI1.XI7.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<11>.MM_i_0_15_63 XI2.XI1.XI7.XI3<11>.DUMMY1 REG_DATA_6<11>
+ XI2.XI1.XI7.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<11>.NEN
+ XI2.XI1.XI7.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<11>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<11>.MM_i_24 VDD! XI2.XI1.XI7.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<11>.MM_i_24_1 XI2.XI1.XI7.XI3<11>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<11>.MM_i_24_0 VDD! REG_DATA_6<11> XI2.XI1.XI7.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI7.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_6<11> XI2.XI1.XI7.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<11>.MM_i_24_1_48 XI2.XI1.XI7.XI3<11>.Y XI2.XI1.XI7.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<11>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<10>.MM_i_0 VSS! XI2.XI1.XI7.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<10>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<10>.MM_i_0_15 VSS! REG_DATA_6<10> XI2.XI1.XI7.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<10>.MM_i_0_15_63 XI2.XI1.XI7.XI3<10>.DUMMY1 REG_DATA_6<10>
+ XI2.XI1.XI7.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<10>.NEN
+ XI2.XI1.XI7.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<10>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<10>.MM_i_24 VDD! XI2.XI1.XI7.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<10>.MM_i_24_1 XI2.XI1.XI7.XI3<10>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<10>.MM_i_24_0 VDD! REG_DATA_6<10> XI2.XI1.XI7.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI7.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_6<10> XI2.XI1.XI7.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<10>.MM_i_24_1_48 XI2.XI1.XI7.XI3<10>.Y XI2.XI1.XI7.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<10>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<9>.MM_i_0 VSS! XI2.XI1.XI7.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<9>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<9>.MM_i_0_15 VSS! REG_DATA_6<9> XI2.XI1.XI7.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<9>.MM_i_0_15_63 XI2.XI1.XI7.XI3<9>.DUMMY1 REG_DATA_6<9>
+ XI2.XI1.XI7.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<9>.NEN
+ XI2.XI1.XI7.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<9>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<9>.MM_i_24 VDD! XI2.XI1.XI7.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<9>.MM_i_24_1 XI2.XI1.XI7.XI3<9>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<9>.MM_i_24_0 VDD! REG_DATA_6<9> XI2.XI1.XI7.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_6<9> XI2.XI1.XI7.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<9>.MM_i_24_1_48 XI2.XI1.XI7.XI3<9>.Y XI2.XI1.XI7.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<9>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<8>.MM_i_0 VSS! XI2.XI1.XI7.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<8>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<8>.MM_i_0_15 VSS! REG_DATA_6<8> XI2.XI1.XI7.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<8>.MM_i_0_15_63 XI2.XI1.XI7.XI3<8>.DUMMY1 REG_DATA_6<8>
+ XI2.XI1.XI7.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<8>.NEN
+ XI2.XI1.XI7.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<8>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<8>.MM_i_24 VDD! XI2.XI1.XI7.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<8>.MM_i_24_1 XI2.XI1.XI7.XI3<8>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<8>.MM_i_24_0 VDD! REG_DATA_6<8> XI2.XI1.XI7.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_6<8> XI2.XI1.XI7.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<8>.MM_i_24_1_48 XI2.XI1.XI7.XI3<8>.Y XI2.XI1.XI7.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<8>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<15>.MM_i_0 VSS! XI2.XI1.XI7.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<15>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<15>.MM_i_0_15 VSS! REG_DATA_6<15> XI2.XI1.XI7.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<15>.MM_i_0_15_63 XI2.XI1.XI7.XI3<15>.DUMMY1 REG_DATA_6<15>
+ XI2.XI1.XI7.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<15>.NEN
+ XI2.XI1.XI7.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<15>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<15>.MM_i_24 VDD! XI2.XI1.XI7.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<15>.MM_i_24_1 XI2.XI1.XI7.XI3<15>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<15>.MM_i_24_0 VDD! REG_DATA_6<15> XI2.XI1.XI7.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI7.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_6<15> XI2.XI1.XI7.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<15>.MM_i_24_1_48 XI2.XI1.XI7.XI3<15>.Y XI2.XI1.XI7.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<15>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<14>.MM_i_0 VSS! XI2.XI1.XI7.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<14>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<14>.MM_i_0_15 VSS! REG_DATA_6<14> XI2.XI1.XI7.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<14>.MM_i_0_15_63 XI2.XI1.XI7.XI3<14>.DUMMY1 REG_DATA_6<14>
+ XI2.XI1.XI7.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<14>.NEN
+ XI2.XI1.XI7.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<14>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<14>.MM_i_24 VDD! XI2.XI1.XI7.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<14>.MM_i_24_1 XI2.XI1.XI7.XI3<14>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<14>.MM_i_24_0 VDD! REG_DATA_6<14> XI2.XI1.XI7.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI7.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_6<14> XI2.XI1.XI7.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<14>.MM_i_24_1_48 XI2.XI1.XI7.XI3<14>.Y XI2.XI1.XI7.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<14>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<13>.MM_i_0 VSS! XI2.XI1.XI7.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<13>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<13>.MM_i_0_15 VSS! REG_DATA_6<13> XI2.XI1.XI7.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<13>.MM_i_0_15_63 XI2.XI1.XI7.XI3<13>.DUMMY1 REG_DATA_6<13>
+ XI2.XI1.XI7.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<13>.NEN
+ XI2.XI1.XI7.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<13>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<13>.MM_i_24 VDD! XI2.XI1.XI7.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<13>.MM_i_24_1 XI2.XI1.XI7.XI3<13>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<13>.MM_i_24_0 VDD! REG_DATA_6<13> XI2.XI1.XI7.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI7.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_6<13> XI2.XI1.XI7.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<13>.MM_i_24_1_48 XI2.XI1.XI7.XI3<13>.Y XI2.XI1.XI7.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<13>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI7.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI7.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI7.XI3<12>.MM_i_0 VSS! XI2.XI1.XI7.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI7.XI3<12>.MM_i_0_14 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<12>.MM_i_0_15 VSS! REG_DATA_6<12> XI2.XI1.XI7.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<12>.MM_i_0_15_63 XI2.XI1.XI7.XI3<12>.DUMMY1 REG_DATA_6<12>
+ XI2.XI1.XI7.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI7.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI7.XI3<12>.NEN
+ XI2.XI1.XI7.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI7.XI3<12>.MM_i_17 VSS! XI2.NET1<6> XI2.XI1.XI7.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI7.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI7.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<12>.MM_i_24 VDD! XI2.XI1.XI7.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI7.XI3<12>.MM_i_24_1 XI2.XI1.XI7.XI3<12>.DUMMY0 XI2.NET1<6>
+ XI2.XI1.XI7.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI7.XI3<12>.MM_i_24_0 VDD! REG_DATA_6<12> XI2.XI1.XI7.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI7.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_6<12> XI2.XI1.XI7.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI7.XI3<12>.MM_i_24_1_48 XI2.XI1.XI7.XI3<12>.Y XI2.XI1.XI7.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI7.XI3<12>.MM_i_42 VDD! XI2.NET1<6> XI2.XI1.XI7.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<3>.MM_i_0 VSS! XI2.XI1.XI8.XI3<3>.X RD_DATA_1<3> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<3>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<3>.MM_i_0_15 VSS! REG_DATA_5<3> XI2.XI1.XI8.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<3>.MM_i_0_15_63 XI2.XI1.XI8.XI3<3>.DUMMY1 REG_DATA_5<3>
+ XI2.XI1.XI8.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<3>.NEN
+ XI2.XI1.XI8.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<3>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<3>.MM_i_24 VDD! XI2.XI1.XI8.XI3<3>.Y RD_DATA_1<3> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<3>.MM_i_24_1 XI2.XI1.XI8.XI3<3>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<3>.MM_i_24_0 VDD! REG_DATA_5<3> XI2.XI1.XI8.XI3<3>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_5<3> XI2.XI1.XI8.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<3>.MM_i_24_1_48 XI2.XI1.XI8.XI3<3>.Y XI2.XI1.XI8.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<3>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<2>.MM_i_0 VSS! XI2.XI1.XI8.XI3<2>.X RD_DATA_1<2> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<2>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<2>.MM_i_0_15 VSS! REG_DATA_5<2> XI2.XI1.XI8.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<2>.MM_i_0_15_63 XI2.XI1.XI8.XI3<2>.DUMMY1 REG_DATA_5<2>
+ XI2.XI1.XI8.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<2>.NEN
+ XI2.XI1.XI8.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<2>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<2>.MM_i_24 VDD! XI2.XI1.XI8.XI3<2>.Y RD_DATA_1<2> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<2>.MM_i_24_1 XI2.XI1.XI8.XI3<2>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<2>.MM_i_24_0 VDD! REG_DATA_5<2> XI2.XI1.XI8.XI3<2>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_5<2> XI2.XI1.XI8.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<2>.MM_i_24_1_48 XI2.XI1.XI8.XI3<2>.Y XI2.XI1.XI8.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<2>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<1>.MM_i_0 VSS! XI2.XI1.XI8.XI3<1>.X RD_DATA_1<1> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<1>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<1>.MM_i_0_15 VSS! REG_DATA_5<1> XI2.XI1.XI8.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<1>.MM_i_0_15_63 XI2.XI1.XI8.XI3<1>.DUMMY1 REG_DATA_5<1>
+ XI2.XI1.XI8.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<1>.NEN
+ XI2.XI1.XI8.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<1>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<1>.MM_i_24 VDD! XI2.XI1.XI8.XI3<1>.Y RD_DATA_1<1> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<1>.MM_i_24_1 XI2.XI1.XI8.XI3<1>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<1>.MM_i_24_0 VDD! REG_DATA_5<1> XI2.XI1.XI8.XI3<1>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_5<1> XI2.XI1.XI8.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<1>.MM_i_24_1_48 XI2.XI1.XI8.XI3<1>.Y XI2.XI1.XI8.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<1>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<0>.MM_i_0 VSS! XI2.XI1.XI8.XI3<0>.X RD_DATA_1<0> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<0>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<0>.MM_i_0_15 VSS! REG_DATA_5<0> XI2.XI1.XI8.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<0>.MM_i_0_15_63 XI2.XI1.XI8.XI3<0>.DUMMY1 REG_DATA_5<0>
+ XI2.XI1.XI8.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<0>.NEN
+ XI2.XI1.XI8.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<0>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<0>.MM_i_24 VDD! XI2.XI1.XI8.XI3<0>.Y RD_DATA_1<0> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<0>.MM_i_24_1 XI2.XI1.XI8.XI3<0>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<0>.MM_i_24_0 VDD! REG_DATA_5<0> XI2.XI1.XI8.XI3<0>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_5<0> XI2.XI1.XI8.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<0>.MM_i_24_1_48 XI2.XI1.XI8.XI3<0>.Y XI2.XI1.XI8.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<0>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<7>.MM_i_0 VSS! XI2.XI1.XI8.XI3<7>.X RD_DATA_1<7> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<7>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<7>.MM_i_0_15 VSS! REG_DATA_5<7> XI2.XI1.XI8.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<7>.MM_i_0_15_63 XI2.XI1.XI8.XI3<7>.DUMMY1 REG_DATA_5<7>
+ XI2.XI1.XI8.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<7>.NEN
+ XI2.XI1.XI8.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<7>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<7>.MM_i_24 VDD! XI2.XI1.XI8.XI3<7>.Y RD_DATA_1<7> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<7>.MM_i_24_1 XI2.XI1.XI8.XI3<7>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<7>.MM_i_24_0 VDD! REG_DATA_5<7> XI2.XI1.XI8.XI3<7>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_5<7> XI2.XI1.XI8.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<7>.MM_i_24_1_48 XI2.XI1.XI8.XI3<7>.Y XI2.XI1.XI8.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<7>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<6>.MM_i_0 VSS! XI2.XI1.XI8.XI3<6>.X RD_DATA_1<6> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<6>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<6>.MM_i_0_15 VSS! REG_DATA_5<6> XI2.XI1.XI8.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<6>.MM_i_0_15_63 XI2.XI1.XI8.XI3<6>.DUMMY1 REG_DATA_5<6>
+ XI2.XI1.XI8.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<6>.NEN
+ XI2.XI1.XI8.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<6>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<6>.MM_i_24 VDD! XI2.XI1.XI8.XI3<6>.Y RD_DATA_1<6> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<6>.MM_i_24_1 XI2.XI1.XI8.XI3<6>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<6>.MM_i_24_0 VDD! REG_DATA_5<6> XI2.XI1.XI8.XI3<6>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_5<6> XI2.XI1.XI8.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<6>.MM_i_24_1_48 XI2.XI1.XI8.XI3<6>.Y XI2.XI1.XI8.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<6>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<5>.MM_i_0 VSS! XI2.XI1.XI8.XI3<5>.X RD_DATA_1<5> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<5>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<5>.MM_i_0_15 VSS! REG_DATA_5<5> XI2.XI1.XI8.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<5>.MM_i_0_15_63 XI2.XI1.XI8.XI3<5>.DUMMY1 REG_DATA_5<5>
+ XI2.XI1.XI8.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<5>.NEN
+ XI2.XI1.XI8.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<5>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<5>.MM_i_24 VDD! XI2.XI1.XI8.XI3<5>.Y RD_DATA_1<5> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<5>.MM_i_24_1 XI2.XI1.XI8.XI3<5>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<5>.MM_i_24_0 VDD! REG_DATA_5<5> XI2.XI1.XI8.XI3<5>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_5<5> XI2.XI1.XI8.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<5>.MM_i_24_1_48 XI2.XI1.XI8.XI3<5>.Y XI2.XI1.XI8.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<5>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<4>.MM_i_0 VSS! XI2.XI1.XI8.XI3<4>.X RD_DATA_1<4> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<4>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<4>.MM_i_0_15 VSS! REG_DATA_5<4> XI2.XI1.XI8.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<4>.MM_i_0_15_63 XI2.XI1.XI8.XI3<4>.DUMMY1 REG_DATA_5<4>
+ XI2.XI1.XI8.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<4>.NEN
+ XI2.XI1.XI8.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<4>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<4>.MM_i_24 VDD! XI2.XI1.XI8.XI3<4>.Y RD_DATA_1<4> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<4>.MM_i_24_1 XI2.XI1.XI8.XI3<4>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<4>.MM_i_24_0 VDD! REG_DATA_5<4> XI2.XI1.XI8.XI3<4>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_5<4> XI2.XI1.XI8.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<4>.MM_i_24_1_48 XI2.XI1.XI8.XI3<4>.Y XI2.XI1.XI8.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<4>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<11>.MM_i_0 VSS! XI2.XI1.XI8.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<11>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<11>.MM_i_0_15 VSS! REG_DATA_5<11> XI2.XI1.XI8.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<11>.MM_i_0_15_63 XI2.XI1.XI8.XI3<11>.DUMMY1 REG_DATA_5<11>
+ XI2.XI1.XI8.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<11>.NEN
+ XI2.XI1.XI8.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<11>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<11>.MM_i_24 VDD! XI2.XI1.XI8.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<11>.MM_i_24_1 XI2.XI1.XI8.XI3<11>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<11>.MM_i_24_0 VDD! REG_DATA_5<11> XI2.XI1.XI8.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI8.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_5<11> XI2.XI1.XI8.XI3<11>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<11>.MM_i_24_1_48 XI2.XI1.XI8.XI3<11>.Y XI2.XI1.XI8.XI3<11>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<11>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<10>.MM_i_0 VSS! XI2.XI1.XI8.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<10>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<10>.MM_i_0_15 VSS! REG_DATA_5<10> XI2.XI1.XI8.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<10>.MM_i_0_15_63 XI2.XI1.XI8.XI3<10>.DUMMY1 REG_DATA_5<10>
+ XI2.XI1.XI8.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<10>.NEN
+ XI2.XI1.XI8.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<10>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<10>.MM_i_24 VDD! XI2.XI1.XI8.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<10>.MM_i_24_1 XI2.XI1.XI8.XI3<10>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<10>.MM_i_24_0 VDD! REG_DATA_5<10> XI2.XI1.XI8.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI8.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_5<10> XI2.XI1.XI8.XI3<10>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<10>.MM_i_24_1_48 XI2.XI1.XI8.XI3<10>.Y XI2.XI1.XI8.XI3<10>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<10>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<9>.MM_i_0 VSS! XI2.XI1.XI8.XI3<9>.X RD_DATA_1<9> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<9>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<9>.MM_i_0_15 VSS! REG_DATA_5<9> XI2.XI1.XI8.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<9>.MM_i_0_15_63 XI2.XI1.XI8.XI3<9>.DUMMY1 REG_DATA_5<9>
+ XI2.XI1.XI8.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<9>.NEN
+ XI2.XI1.XI8.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<9>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<9>.MM_i_24 VDD! XI2.XI1.XI8.XI3<9>.Y RD_DATA_1<9> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<9>.MM_i_24_1 XI2.XI1.XI8.XI3<9>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<9>.MM_i_24_0 VDD! REG_DATA_5<9> XI2.XI1.XI8.XI3<9>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_5<9> XI2.XI1.XI8.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<9>.MM_i_24_1_48 XI2.XI1.XI8.XI3<9>.Y XI2.XI1.XI8.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<9>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<8>.MM_i_0 VSS! XI2.XI1.XI8.XI3<8>.X RD_DATA_1<8> VSS! NMOS_VTL
+ L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<8>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<8>.MM_i_0_15 VSS! REG_DATA_5<8> XI2.XI1.XI8.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<8>.MM_i_0_15_63 XI2.XI1.XI8.XI3<8>.DUMMY1 REG_DATA_5<8>
+ XI2.XI1.XI8.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<8>.NEN
+ XI2.XI1.XI8.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<8>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<8>.MM_i_24 VDD! XI2.XI1.XI8.XI3<8>.Y RD_DATA_1<8> VDD! PMOS_VTL
+ L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<8>.MM_i_24_1 XI2.XI1.XI8.XI3<8>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<8>.MM_i_24_0 VDD! REG_DATA_5<8> XI2.XI1.XI8.XI3<8>.DUMMY0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_5<8> XI2.XI1.XI8.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<8>.MM_i_24_1_48 XI2.XI1.XI8.XI3<8>.Y XI2.XI1.XI8.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<8>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<15>.MM_i_0 VSS! XI2.XI1.XI8.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<15>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<15>.MM_i_0_15 VSS! REG_DATA_5<15> XI2.XI1.XI8.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<15>.MM_i_0_15_63 XI2.XI1.XI8.XI3<15>.DUMMY1 REG_DATA_5<15>
+ XI2.XI1.XI8.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<15>.NEN
+ XI2.XI1.XI8.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<15>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<15>.MM_i_24 VDD! XI2.XI1.XI8.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<15>.MM_i_24_1 XI2.XI1.XI8.XI3<15>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<15>.MM_i_24_0 VDD! REG_DATA_5<15> XI2.XI1.XI8.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI8.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_5<15> XI2.XI1.XI8.XI3<15>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<15>.MM_i_24_1_48 XI2.XI1.XI8.XI3<15>.Y XI2.XI1.XI8.XI3<15>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<15>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<14>.MM_i_0 VSS! XI2.XI1.XI8.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<14>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<14>.MM_i_0_15 VSS! REG_DATA_5<14> XI2.XI1.XI8.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<14>.MM_i_0_15_63 XI2.XI1.XI8.XI3<14>.DUMMY1 REG_DATA_5<14>
+ XI2.XI1.XI8.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<14>.NEN
+ XI2.XI1.XI8.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<14>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<14>.MM_i_24 VDD! XI2.XI1.XI8.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<14>.MM_i_24_1 XI2.XI1.XI8.XI3<14>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<14>.MM_i_24_0 VDD! REG_DATA_5<14> XI2.XI1.XI8.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI8.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_5<14> XI2.XI1.XI8.XI3<14>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<14>.MM_i_24_1_48 XI2.XI1.XI8.XI3<14>.Y XI2.XI1.XI8.XI3<14>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<14>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<13>.MM_i_0 VSS! XI2.XI1.XI8.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<13>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<13>.MM_i_0_15 VSS! REG_DATA_5<13> XI2.XI1.XI8.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<13>.MM_i_0_15_63 XI2.XI1.XI8.XI3<13>.DUMMY1 REG_DATA_5<13>
+ XI2.XI1.XI8.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<13>.NEN
+ XI2.XI1.XI8.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<13>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<13>.MM_i_24 VDD! XI2.XI1.XI8.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<13>.MM_i_24_1 XI2.XI1.XI8.XI3<13>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<13>.MM_i_24_0 VDD! REG_DATA_5<13> XI2.XI1.XI8.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI8.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_5<13> XI2.XI1.XI8.XI3<13>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<13>.MM_i_24_1_48 XI2.XI1.XI8.XI3<13>.Y XI2.XI1.XI8.XI3<13>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<13>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI8.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI8.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI8.XI3<12>.MM_i_0 VSS! XI2.XI1.XI8.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI8.XI3<12>.MM_i_0_14 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<12>.MM_i_0_15 VSS! REG_DATA_5<12> XI2.XI1.XI8.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<12>.MM_i_0_15_63 XI2.XI1.XI8.XI3<12>.DUMMY1 REG_DATA_5<12>
+ XI2.XI1.XI8.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI8.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI8.XI3<12>.NEN
+ XI2.XI1.XI8.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI8.XI3<12>.MM_i_17 VSS! XI2.NET1<7> XI2.XI1.XI8.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI8.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI8.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<12>.MM_i_24 VDD! XI2.XI1.XI8.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI8.XI3<12>.MM_i_24_1 XI2.XI1.XI8.XI3<12>.DUMMY0 XI2.NET1<7>
+ XI2.XI1.XI8.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI8.XI3<12>.MM_i_24_0 VDD! REG_DATA_5<12> XI2.XI1.XI8.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI8.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_5<12> XI2.XI1.XI8.XI3<12>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI8.XI3<12>.MM_i_24_1_48 XI2.XI1.XI8.XI3<12>.Y XI2.XI1.XI8.XI3<12>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI8.XI3<12>.MM_i_42 VDD! XI2.NET1<7> XI2.XI1.XI8.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<3>.MM_i_0 VSS! XI2.XI1.XI11.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<3>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<3>.MM_i_0_15 VSS! REG_DATA_4<3> XI2.XI1.XI11.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<3>.MM_i_0_15_63 XI2.XI1.XI11.XI3<3>.DUMMY1 REG_DATA_4<3>
+ XI2.XI1.XI11.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<3>.NEN
+ XI2.XI1.XI11.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<3>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<3>.MM_i_24 VDD! XI2.XI1.XI11.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<3>.MM_i_24_1 XI2.XI1.XI11.XI3<3>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<3>.MM_i_24_0 VDD! REG_DATA_4<3> XI2.XI1.XI11.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_4<3> XI2.XI1.XI11.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<3>.MM_i_24_1_48 XI2.XI1.XI11.XI3<3>.Y XI2.XI1.XI11.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<3>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<2>.MM_i_0 VSS! XI2.XI1.XI11.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<2>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<2>.MM_i_0_15 VSS! REG_DATA_4<2> XI2.XI1.XI11.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<2>.MM_i_0_15_63 XI2.XI1.XI11.XI3<2>.DUMMY1 REG_DATA_4<2>
+ XI2.XI1.XI11.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<2>.NEN
+ XI2.XI1.XI11.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<2>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<2>.MM_i_24 VDD! XI2.XI1.XI11.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<2>.MM_i_24_1 XI2.XI1.XI11.XI3<2>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<2>.MM_i_24_0 VDD! REG_DATA_4<2> XI2.XI1.XI11.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_4<2> XI2.XI1.XI11.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<2>.MM_i_24_1_48 XI2.XI1.XI11.XI3<2>.Y XI2.XI1.XI11.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<2>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<1>.MM_i_0 VSS! XI2.XI1.XI11.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<1>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<1>.MM_i_0_15 VSS! REG_DATA_4<1> XI2.XI1.XI11.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<1>.MM_i_0_15_63 XI2.XI1.XI11.XI3<1>.DUMMY1 REG_DATA_4<1>
+ XI2.XI1.XI11.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<1>.NEN
+ XI2.XI1.XI11.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<1>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<1>.MM_i_24 VDD! XI2.XI1.XI11.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<1>.MM_i_24_1 XI2.XI1.XI11.XI3<1>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<1>.MM_i_24_0 VDD! REG_DATA_4<1> XI2.XI1.XI11.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_4<1> XI2.XI1.XI11.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<1>.MM_i_24_1_48 XI2.XI1.XI11.XI3<1>.Y XI2.XI1.XI11.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<1>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<0>.MM_i_0 VSS! XI2.XI1.XI11.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<0>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<0>.MM_i_0_15 VSS! REG_DATA_4<0> XI2.XI1.XI11.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<0>.MM_i_0_15_63 XI2.XI1.XI11.XI3<0>.DUMMY1 REG_DATA_4<0>
+ XI2.XI1.XI11.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<0>.NEN
+ XI2.XI1.XI11.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<0>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<0>.MM_i_24 VDD! XI2.XI1.XI11.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<0>.MM_i_24_1 XI2.XI1.XI11.XI3<0>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<0>.MM_i_24_0 VDD! REG_DATA_4<0> XI2.XI1.XI11.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_4<0> XI2.XI1.XI11.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<0>.MM_i_24_1_48 XI2.XI1.XI11.XI3<0>.Y XI2.XI1.XI11.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<0>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<7>.MM_i_0 VSS! XI2.XI1.XI11.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<7>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<7>.MM_i_0_15 VSS! REG_DATA_4<7> XI2.XI1.XI11.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<7>.MM_i_0_15_63 XI2.XI1.XI11.XI3<7>.DUMMY1 REG_DATA_4<7>
+ XI2.XI1.XI11.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<7>.NEN
+ XI2.XI1.XI11.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<7>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<7>.MM_i_24 VDD! XI2.XI1.XI11.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<7>.MM_i_24_1 XI2.XI1.XI11.XI3<7>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<7>.MM_i_24_0 VDD! REG_DATA_4<7> XI2.XI1.XI11.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_4<7> XI2.XI1.XI11.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<7>.MM_i_24_1_48 XI2.XI1.XI11.XI3<7>.Y XI2.XI1.XI11.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<7>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<6>.MM_i_0 VSS! XI2.XI1.XI11.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<6>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<6>.MM_i_0_15 VSS! REG_DATA_4<6> XI2.XI1.XI11.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<6>.MM_i_0_15_63 XI2.XI1.XI11.XI3<6>.DUMMY1 REG_DATA_4<6>
+ XI2.XI1.XI11.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<6>.NEN
+ XI2.XI1.XI11.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<6>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<6>.MM_i_24 VDD! XI2.XI1.XI11.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<6>.MM_i_24_1 XI2.XI1.XI11.XI3<6>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<6>.MM_i_24_0 VDD! REG_DATA_4<6> XI2.XI1.XI11.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_4<6> XI2.XI1.XI11.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<6>.MM_i_24_1_48 XI2.XI1.XI11.XI3<6>.Y XI2.XI1.XI11.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<6>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<5>.MM_i_0 VSS! XI2.XI1.XI11.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<5>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<5>.MM_i_0_15 VSS! REG_DATA_4<5> XI2.XI1.XI11.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<5>.MM_i_0_15_63 XI2.XI1.XI11.XI3<5>.DUMMY1 REG_DATA_4<5>
+ XI2.XI1.XI11.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<5>.NEN
+ XI2.XI1.XI11.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<5>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<5>.MM_i_24 VDD! XI2.XI1.XI11.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<5>.MM_i_24_1 XI2.XI1.XI11.XI3<5>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<5>.MM_i_24_0 VDD! REG_DATA_4<5> XI2.XI1.XI11.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_4<5> XI2.XI1.XI11.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<5>.MM_i_24_1_48 XI2.XI1.XI11.XI3<5>.Y XI2.XI1.XI11.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<5>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<4>.MM_i_0 VSS! XI2.XI1.XI11.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<4>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<4>.MM_i_0_15 VSS! REG_DATA_4<4> XI2.XI1.XI11.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<4>.MM_i_0_15_63 XI2.XI1.XI11.XI3<4>.DUMMY1 REG_DATA_4<4>
+ XI2.XI1.XI11.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<4>.NEN
+ XI2.XI1.XI11.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<4>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<4>.MM_i_24 VDD! XI2.XI1.XI11.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<4>.MM_i_24_1 XI2.XI1.XI11.XI3<4>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<4>.MM_i_24_0 VDD! REG_DATA_4<4> XI2.XI1.XI11.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_4<4> XI2.XI1.XI11.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<4>.MM_i_24_1_48 XI2.XI1.XI11.XI3<4>.Y XI2.XI1.XI11.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<4>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<11>.MM_i_0 VSS! XI2.XI1.XI11.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<11>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<11>.MM_i_0_15 VSS! REG_DATA_4<11> XI2.XI1.XI11.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<11>.MM_i_0_15_63 XI2.XI1.XI11.XI3<11>.DUMMY1 REG_DATA_4<11>
+ XI2.XI1.XI11.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<11>.NEN
+ XI2.XI1.XI11.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<11>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<11>.MM_i_24 VDD! XI2.XI1.XI11.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<11>.MM_i_24_1 XI2.XI1.XI11.XI3<11>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<11>.MM_i_24_0 VDD! REG_DATA_4<11> XI2.XI1.XI11.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_4<11> XI2.XI1.XI11.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<11>.MM_i_24_1_48 XI2.XI1.XI11.XI3<11>.Y
+ XI2.XI1.XI11.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI11.XI3<11>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<10>.MM_i_0 VSS! XI2.XI1.XI11.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<10>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<10>.MM_i_0_15 VSS! REG_DATA_4<10> XI2.XI1.XI11.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<10>.MM_i_0_15_63 XI2.XI1.XI11.XI3<10>.DUMMY1 REG_DATA_4<10>
+ XI2.XI1.XI11.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<10>.NEN
+ XI2.XI1.XI11.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<10>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<10>.MM_i_24 VDD! XI2.XI1.XI11.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<10>.MM_i_24_1 XI2.XI1.XI11.XI3<10>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<10>.MM_i_24_0 VDD! REG_DATA_4<10> XI2.XI1.XI11.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_4<10> XI2.XI1.XI11.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<10>.MM_i_24_1_48 XI2.XI1.XI11.XI3<10>.Y
+ XI2.XI1.XI11.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI11.XI3<10>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<9>.MM_i_0 VSS! XI2.XI1.XI11.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<9>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<9>.MM_i_0_15 VSS! REG_DATA_4<9> XI2.XI1.XI11.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<9>.MM_i_0_15_63 XI2.XI1.XI11.XI3<9>.DUMMY1 REG_DATA_4<9>
+ XI2.XI1.XI11.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<9>.NEN
+ XI2.XI1.XI11.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<9>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<9>.MM_i_24 VDD! XI2.XI1.XI11.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<9>.MM_i_24_1 XI2.XI1.XI11.XI3<9>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<9>.MM_i_24_0 VDD! REG_DATA_4<9> XI2.XI1.XI11.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_4<9> XI2.XI1.XI11.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<9>.MM_i_24_1_48 XI2.XI1.XI11.XI3<9>.Y XI2.XI1.XI11.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<9>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<8>.MM_i_0 VSS! XI2.XI1.XI11.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<8>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<8>.MM_i_0_15 VSS! REG_DATA_4<8> XI2.XI1.XI11.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<8>.MM_i_0_15_63 XI2.XI1.XI11.XI3<8>.DUMMY1 REG_DATA_4<8>
+ XI2.XI1.XI11.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<8>.NEN
+ XI2.XI1.XI11.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<8>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<8>.MM_i_24 VDD! XI2.XI1.XI11.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<8>.MM_i_24_1 XI2.XI1.XI11.XI3<8>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<8>.MM_i_24_0 VDD! REG_DATA_4<8> XI2.XI1.XI11.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_4<8> XI2.XI1.XI11.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI11.XI3<8>.MM_i_24_1_48 XI2.XI1.XI11.XI3<8>.Y XI2.XI1.XI11.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI11.XI3<8>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<15>.MM_i_0 VSS! XI2.XI1.XI11.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<15>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<15>.MM_i_0_15 VSS! REG_DATA_4<15> XI2.XI1.XI11.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<15>.MM_i_0_15_63 XI2.XI1.XI11.XI3<15>.DUMMY1 REG_DATA_4<15>
+ XI2.XI1.XI11.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<15>.NEN
+ XI2.XI1.XI11.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<15>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<15>.MM_i_24 VDD! XI2.XI1.XI11.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<15>.MM_i_24_1 XI2.XI1.XI11.XI3<15>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<15>.MM_i_24_0 VDD! REG_DATA_4<15> XI2.XI1.XI11.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_4<15> XI2.XI1.XI11.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<15>.MM_i_24_1_48 XI2.XI1.XI11.XI3<15>.Y
+ XI2.XI1.XI11.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI11.XI3<15>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<14>.MM_i_0 VSS! XI2.XI1.XI11.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<14>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<14>.MM_i_0_15 VSS! REG_DATA_4<14> XI2.XI1.XI11.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<14>.MM_i_0_15_63 XI2.XI1.XI11.XI3<14>.DUMMY1 REG_DATA_4<14>
+ XI2.XI1.XI11.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<14>.NEN
+ XI2.XI1.XI11.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<14>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<14>.MM_i_24 VDD! XI2.XI1.XI11.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<14>.MM_i_24_1 XI2.XI1.XI11.XI3<14>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<14>.MM_i_24_0 VDD! REG_DATA_4<14> XI2.XI1.XI11.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_4<14> XI2.XI1.XI11.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<14>.MM_i_24_1_48 XI2.XI1.XI11.XI3<14>.Y
+ XI2.XI1.XI11.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI11.XI3<14>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<13>.MM_i_0 VSS! XI2.XI1.XI11.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<13>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<13>.MM_i_0_15 VSS! REG_DATA_4<13> XI2.XI1.XI11.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<13>.MM_i_0_15_63 XI2.XI1.XI11.XI3<13>.DUMMY1 REG_DATA_4<13>
+ XI2.XI1.XI11.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<13>.NEN
+ XI2.XI1.XI11.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<13>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<13>.MM_i_24 VDD! XI2.XI1.XI11.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<13>.MM_i_24_1 XI2.XI1.XI11.XI3<13>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<13>.MM_i_24_0 VDD! REG_DATA_4<13> XI2.XI1.XI11.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_4<13> XI2.XI1.XI11.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<13>.MM_i_24_1_48 XI2.XI1.XI11.XI3<13>.Y
+ XI2.XI1.XI11.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI11.XI3<13>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI11.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI11.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI11.XI3<12>.MM_i_0 VSS! XI2.XI1.XI11.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI11.XI3<12>.MM_i_0_14 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<12>.MM_i_0_15 VSS! REG_DATA_4<12> XI2.XI1.XI11.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<12>.MM_i_0_15_63 XI2.XI1.XI11.XI3<12>.DUMMY1 REG_DATA_4<12>
+ XI2.XI1.XI11.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI11.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI11.XI3<12>.NEN
+ XI2.XI1.XI11.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI11.XI3<12>.MM_i_17 VSS! XI2.NET1<8> XI2.XI1.XI11.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI11.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI11.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<12>.MM_i_24 VDD! XI2.XI1.XI11.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI11.XI3<12>.MM_i_24_1 XI2.XI1.XI11.XI3<12>.DUMMY0 XI2.NET1<8>
+ XI2.XI1.XI11.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI11.XI3<12>.MM_i_24_0 VDD! REG_DATA_4<12> XI2.XI1.XI11.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_4<12> XI2.XI1.XI11.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI11.XI3<12>.MM_i_24_1_48 XI2.XI1.XI11.XI3<12>.Y
+ XI2.XI1.XI11.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI11.XI3<12>.MM_i_42 VDD! XI2.NET1<8> XI2.XI1.XI11.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<3>.MM_i_0 VSS! XI2.XI1.XI12.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<3>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<3>.MM_i_0_15 VSS! REG_DATA_3<3> XI2.XI1.XI12.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<3>.MM_i_0_15_63 XI2.XI1.XI12.XI3<3>.DUMMY1 REG_DATA_3<3>
+ XI2.XI1.XI12.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<3>.NEN
+ XI2.XI1.XI12.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<3>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<3>.MM_i_24 VDD! XI2.XI1.XI12.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<3>.MM_i_24_1 XI2.XI1.XI12.XI3<3>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<3>.MM_i_24_0 VDD! REG_DATA_3<3> XI2.XI1.XI12.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_3<3> XI2.XI1.XI12.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<3>.MM_i_24_1_48 XI2.XI1.XI12.XI3<3>.Y XI2.XI1.XI12.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<3>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<2>.MM_i_0 VSS! XI2.XI1.XI12.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<2>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<2>.MM_i_0_15 VSS! REG_DATA_3<2> XI2.XI1.XI12.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<2>.MM_i_0_15_63 XI2.XI1.XI12.XI3<2>.DUMMY1 REG_DATA_3<2>
+ XI2.XI1.XI12.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<2>.NEN
+ XI2.XI1.XI12.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<2>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<2>.MM_i_24 VDD! XI2.XI1.XI12.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<2>.MM_i_24_1 XI2.XI1.XI12.XI3<2>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<2>.MM_i_24_0 VDD! REG_DATA_3<2> XI2.XI1.XI12.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_3<2> XI2.XI1.XI12.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<2>.MM_i_24_1_48 XI2.XI1.XI12.XI3<2>.Y XI2.XI1.XI12.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<2>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<1>.MM_i_0 VSS! XI2.XI1.XI12.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<1>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<1>.MM_i_0_15 VSS! REG_DATA_3<1> XI2.XI1.XI12.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<1>.MM_i_0_15_63 XI2.XI1.XI12.XI3<1>.DUMMY1 REG_DATA_3<1>
+ XI2.XI1.XI12.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<1>.NEN
+ XI2.XI1.XI12.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<1>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<1>.MM_i_24 VDD! XI2.XI1.XI12.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<1>.MM_i_24_1 XI2.XI1.XI12.XI3<1>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<1>.MM_i_24_0 VDD! REG_DATA_3<1> XI2.XI1.XI12.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_3<1> XI2.XI1.XI12.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<1>.MM_i_24_1_48 XI2.XI1.XI12.XI3<1>.Y XI2.XI1.XI12.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<1>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<0>.MM_i_0 VSS! XI2.XI1.XI12.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<0>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<0>.MM_i_0_15 VSS! REG_DATA_3<0> XI2.XI1.XI12.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<0>.MM_i_0_15_63 XI2.XI1.XI12.XI3<0>.DUMMY1 REG_DATA_3<0>
+ XI2.XI1.XI12.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<0>.NEN
+ XI2.XI1.XI12.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<0>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<0>.MM_i_24 VDD! XI2.XI1.XI12.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<0>.MM_i_24_1 XI2.XI1.XI12.XI3<0>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<0>.MM_i_24_0 VDD! REG_DATA_3<0> XI2.XI1.XI12.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_3<0> XI2.XI1.XI12.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<0>.MM_i_24_1_48 XI2.XI1.XI12.XI3<0>.Y XI2.XI1.XI12.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<0>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<7>.MM_i_0 VSS! XI2.XI1.XI12.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<7>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<7>.MM_i_0_15 VSS! REG_DATA_3<7> XI2.XI1.XI12.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<7>.MM_i_0_15_63 XI2.XI1.XI12.XI3<7>.DUMMY1 REG_DATA_3<7>
+ XI2.XI1.XI12.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<7>.NEN
+ XI2.XI1.XI12.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<7>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<7>.MM_i_24 VDD! XI2.XI1.XI12.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<7>.MM_i_24_1 XI2.XI1.XI12.XI3<7>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<7>.MM_i_24_0 VDD! REG_DATA_3<7> XI2.XI1.XI12.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_3<7> XI2.XI1.XI12.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<7>.MM_i_24_1_48 XI2.XI1.XI12.XI3<7>.Y XI2.XI1.XI12.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<7>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<6>.MM_i_0 VSS! XI2.XI1.XI12.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<6>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<6>.MM_i_0_15 VSS! REG_DATA_3<6> XI2.XI1.XI12.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<6>.MM_i_0_15_63 XI2.XI1.XI12.XI3<6>.DUMMY1 REG_DATA_3<6>
+ XI2.XI1.XI12.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<6>.NEN
+ XI2.XI1.XI12.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<6>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<6>.MM_i_24 VDD! XI2.XI1.XI12.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<6>.MM_i_24_1 XI2.XI1.XI12.XI3<6>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<6>.MM_i_24_0 VDD! REG_DATA_3<6> XI2.XI1.XI12.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_3<6> XI2.XI1.XI12.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<6>.MM_i_24_1_48 XI2.XI1.XI12.XI3<6>.Y XI2.XI1.XI12.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<6>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<5>.MM_i_0 VSS! XI2.XI1.XI12.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<5>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<5>.MM_i_0_15 VSS! REG_DATA_3<5> XI2.XI1.XI12.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<5>.MM_i_0_15_63 XI2.XI1.XI12.XI3<5>.DUMMY1 REG_DATA_3<5>
+ XI2.XI1.XI12.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<5>.NEN
+ XI2.XI1.XI12.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<5>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<5>.MM_i_24 VDD! XI2.XI1.XI12.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<5>.MM_i_24_1 XI2.XI1.XI12.XI3<5>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<5>.MM_i_24_0 VDD! REG_DATA_3<5> XI2.XI1.XI12.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_3<5> XI2.XI1.XI12.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<5>.MM_i_24_1_48 XI2.XI1.XI12.XI3<5>.Y XI2.XI1.XI12.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<5>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<4>.MM_i_0 VSS! XI2.XI1.XI12.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<4>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<4>.MM_i_0_15 VSS! REG_DATA_3<4> XI2.XI1.XI12.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<4>.MM_i_0_15_63 XI2.XI1.XI12.XI3<4>.DUMMY1 REG_DATA_3<4>
+ XI2.XI1.XI12.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<4>.NEN
+ XI2.XI1.XI12.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<4>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<4>.MM_i_24 VDD! XI2.XI1.XI12.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<4>.MM_i_24_1 XI2.XI1.XI12.XI3<4>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<4>.MM_i_24_0 VDD! REG_DATA_3<4> XI2.XI1.XI12.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_3<4> XI2.XI1.XI12.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<4>.MM_i_24_1_48 XI2.XI1.XI12.XI3<4>.Y XI2.XI1.XI12.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<4>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<11>.MM_i_0 VSS! XI2.XI1.XI12.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<11>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<11>.MM_i_0_15 VSS! REG_DATA_3<11> XI2.XI1.XI12.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<11>.MM_i_0_15_63 XI2.XI1.XI12.XI3<11>.DUMMY1 REG_DATA_3<11>
+ XI2.XI1.XI12.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<11>.NEN
+ XI2.XI1.XI12.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<11>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<11>.MM_i_24 VDD! XI2.XI1.XI12.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<11>.MM_i_24_1 XI2.XI1.XI12.XI3<11>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<11>.MM_i_24_0 VDD! REG_DATA_3<11> XI2.XI1.XI12.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_3<11> XI2.XI1.XI12.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<11>.MM_i_24_1_48 XI2.XI1.XI12.XI3<11>.Y
+ XI2.XI1.XI12.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI12.XI3<11>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<10>.MM_i_0 VSS! XI2.XI1.XI12.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<10>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<10>.MM_i_0_15 VSS! REG_DATA_3<10> XI2.XI1.XI12.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<10>.MM_i_0_15_63 XI2.XI1.XI12.XI3<10>.DUMMY1 REG_DATA_3<10>
+ XI2.XI1.XI12.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<10>.NEN
+ XI2.XI1.XI12.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<10>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<10>.MM_i_24 VDD! XI2.XI1.XI12.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<10>.MM_i_24_1 XI2.XI1.XI12.XI3<10>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<10>.MM_i_24_0 VDD! REG_DATA_3<10> XI2.XI1.XI12.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_3<10> XI2.XI1.XI12.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<10>.MM_i_24_1_48 XI2.XI1.XI12.XI3<10>.Y
+ XI2.XI1.XI12.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI12.XI3<10>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<9>.MM_i_0 VSS! XI2.XI1.XI12.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<9>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<9>.MM_i_0_15 VSS! REG_DATA_3<9> XI2.XI1.XI12.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<9>.MM_i_0_15_63 XI2.XI1.XI12.XI3<9>.DUMMY1 REG_DATA_3<9>
+ XI2.XI1.XI12.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<9>.NEN
+ XI2.XI1.XI12.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<9>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<9>.MM_i_24 VDD! XI2.XI1.XI12.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<9>.MM_i_24_1 XI2.XI1.XI12.XI3<9>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<9>.MM_i_24_0 VDD! REG_DATA_3<9> XI2.XI1.XI12.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_3<9> XI2.XI1.XI12.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<9>.MM_i_24_1_48 XI2.XI1.XI12.XI3<9>.Y XI2.XI1.XI12.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<9>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<8>.MM_i_0 VSS! XI2.XI1.XI12.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<8>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<8>.MM_i_0_15 VSS! REG_DATA_3<8> XI2.XI1.XI12.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<8>.MM_i_0_15_63 XI2.XI1.XI12.XI3<8>.DUMMY1 REG_DATA_3<8>
+ XI2.XI1.XI12.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<8>.NEN
+ XI2.XI1.XI12.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<8>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<8>.MM_i_24 VDD! XI2.XI1.XI12.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<8>.MM_i_24_1 XI2.XI1.XI12.XI3<8>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<8>.MM_i_24_0 VDD! REG_DATA_3<8> XI2.XI1.XI12.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_3<8> XI2.XI1.XI12.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI12.XI3<8>.MM_i_24_1_48 XI2.XI1.XI12.XI3<8>.Y XI2.XI1.XI12.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI12.XI3<8>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<15>.MM_i_0 VSS! XI2.XI1.XI12.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<15>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<15>.MM_i_0_15 VSS! REG_DATA_3<15> XI2.XI1.XI12.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<15>.MM_i_0_15_63 XI2.XI1.XI12.XI3<15>.DUMMY1 REG_DATA_3<15>
+ XI2.XI1.XI12.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<15>.NEN
+ XI2.XI1.XI12.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<15>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<15>.MM_i_24 VDD! XI2.XI1.XI12.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<15>.MM_i_24_1 XI2.XI1.XI12.XI3<15>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<15>.MM_i_24_0 VDD! REG_DATA_3<15> XI2.XI1.XI12.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_3<15> XI2.XI1.XI12.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<15>.MM_i_24_1_48 XI2.XI1.XI12.XI3<15>.Y
+ XI2.XI1.XI12.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI12.XI3<15>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<14>.MM_i_0 VSS! XI2.XI1.XI12.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<14>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<14>.MM_i_0_15 VSS! REG_DATA_3<14> XI2.XI1.XI12.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<14>.MM_i_0_15_63 XI2.XI1.XI12.XI3<14>.DUMMY1 REG_DATA_3<14>
+ XI2.XI1.XI12.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<14>.NEN
+ XI2.XI1.XI12.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<14>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<14>.MM_i_24 VDD! XI2.XI1.XI12.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<14>.MM_i_24_1 XI2.XI1.XI12.XI3<14>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<14>.MM_i_24_0 VDD! REG_DATA_3<14> XI2.XI1.XI12.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_3<14> XI2.XI1.XI12.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<14>.MM_i_24_1_48 XI2.XI1.XI12.XI3<14>.Y
+ XI2.XI1.XI12.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI12.XI3<14>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<13>.MM_i_0 VSS! XI2.XI1.XI12.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<13>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<13>.MM_i_0_15 VSS! REG_DATA_3<13> XI2.XI1.XI12.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<13>.MM_i_0_15_63 XI2.XI1.XI12.XI3<13>.DUMMY1 REG_DATA_3<13>
+ XI2.XI1.XI12.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<13>.NEN
+ XI2.XI1.XI12.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<13>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<13>.MM_i_24 VDD! XI2.XI1.XI12.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<13>.MM_i_24_1 XI2.XI1.XI12.XI3<13>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<13>.MM_i_24_0 VDD! REG_DATA_3<13> XI2.XI1.XI12.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_3<13> XI2.XI1.XI12.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<13>.MM_i_24_1_48 XI2.XI1.XI12.XI3<13>.Y
+ XI2.XI1.XI12.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI12.XI3<13>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI12.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI12.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI12.XI3<12>.MM_i_0 VSS! XI2.XI1.XI12.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI12.XI3<12>.MM_i_0_14 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<12>.MM_i_0_15 VSS! REG_DATA_3<12> XI2.XI1.XI12.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<12>.MM_i_0_15_63 XI2.XI1.XI12.XI3<12>.DUMMY1 REG_DATA_3<12>
+ XI2.XI1.XI12.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI12.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI12.XI3<12>.NEN
+ XI2.XI1.XI12.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI12.XI3<12>.MM_i_17 VSS! XI2.NET1<9> XI2.XI1.XI12.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI12.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI12.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<12>.MM_i_24 VDD! XI2.XI1.XI12.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI12.XI3<12>.MM_i_24_1 XI2.XI1.XI12.XI3<12>.DUMMY0 XI2.NET1<9>
+ XI2.XI1.XI12.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI12.XI3<12>.MM_i_24_0 VDD! REG_DATA_3<12> XI2.XI1.XI12.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_3<12> XI2.XI1.XI12.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI12.XI3<12>.MM_i_24_1_48 XI2.XI1.XI12.XI3<12>.Y
+ XI2.XI1.XI12.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI12.XI3<12>.MM_i_42 VDD! XI2.NET1<9> XI2.XI1.XI12.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<3>.MM_i_0 VSS! XI2.XI1.XI14.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<3>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<3>.MM_i_0_15 VSS! REG_DATA_2<3> XI2.XI1.XI14.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<3>.MM_i_0_15_63 XI2.XI1.XI14.XI3<3>.DUMMY1 REG_DATA_2<3>
+ XI2.XI1.XI14.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<3>.NEN
+ XI2.XI1.XI14.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<3>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<3>.MM_i_24 VDD! XI2.XI1.XI14.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<3>.MM_i_24_1 XI2.XI1.XI14.XI3<3>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<3>.MM_i_24_0 VDD! REG_DATA_2<3> XI2.XI1.XI14.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_2<3> XI2.XI1.XI14.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<3>.MM_i_24_1_48 XI2.XI1.XI14.XI3<3>.Y XI2.XI1.XI14.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<3>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<2>.MM_i_0 VSS! XI2.XI1.XI14.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<2>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<2>.MM_i_0_15 VSS! REG_DATA_2<2> XI2.XI1.XI14.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<2>.MM_i_0_15_63 XI2.XI1.XI14.XI3<2>.DUMMY1 REG_DATA_2<2>
+ XI2.XI1.XI14.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<2>.NEN
+ XI2.XI1.XI14.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<2>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<2>.MM_i_24 VDD! XI2.XI1.XI14.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<2>.MM_i_24_1 XI2.XI1.XI14.XI3<2>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<2>.MM_i_24_0 VDD! REG_DATA_2<2> XI2.XI1.XI14.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_2<2> XI2.XI1.XI14.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<2>.MM_i_24_1_48 XI2.XI1.XI14.XI3<2>.Y XI2.XI1.XI14.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<2>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<1>.MM_i_0 VSS! XI2.XI1.XI14.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<1>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<1>.MM_i_0_15 VSS! REG_DATA_2<1> XI2.XI1.XI14.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<1>.MM_i_0_15_63 XI2.XI1.XI14.XI3<1>.DUMMY1 REG_DATA_2<1>
+ XI2.XI1.XI14.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<1>.NEN
+ XI2.XI1.XI14.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<1>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<1>.MM_i_24 VDD! XI2.XI1.XI14.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<1>.MM_i_24_1 XI2.XI1.XI14.XI3<1>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<1>.MM_i_24_0 VDD! REG_DATA_2<1> XI2.XI1.XI14.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_2<1> XI2.XI1.XI14.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<1>.MM_i_24_1_48 XI2.XI1.XI14.XI3<1>.Y XI2.XI1.XI14.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<1>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<0>.MM_i_0 VSS! XI2.XI1.XI14.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<0>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<0>.MM_i_0_15 VSS! REG_DATA_2<0> XI2.XI1.XI14.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<0>.MM_i_0_15_63 XI2.XI1.XI14.XI3<0>.DUMMY1 REG_DATA_2<0>
+ XI2.XI1.XI14.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<0>.NEN
+ XI2.XI1.XI14.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<0>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<0>.MM_i_24 VDD! XI2.XI1.XI14.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<0>.MM_i_24_1 XI2.XI1.XI14.XI3<0>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<0>.MM_i_24_0 VDD! REG_DATA_2<0> XI2.XI1.XI14.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_2<0> XI2.XI1.XI14.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<0>.MM_i_24_1_48 XI2.XI1.XI14.XI3<0>.Y XI2.XI1.XI14.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<0>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<7>.MM_i_0 VSS! XI2.XI1.XI14.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<7>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<7>.MM_i_0_15 VSS! REG_DATA_2<7> XI2.XI1.XI14.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<7>.MM_i_0_15_63 XI2.XI1.XI14.XI3<7>.DUMMY1 REG_DATA_2<7>
+ XI2.XI1.XI14.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<7>.NEN
+ XI2.XI1.XI14.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<7>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<7>.MM_i_24 VDD! XI2.XI1.XI14.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<7>.MM_i_24_1 XI2.XI1.XI14.XI3<7>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<7>.MM_i_24_0 VDD! REG_DATA_2<7> XI2.XI1.XI14.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_2<7> XI2.XI1.XI14.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<7>.MM_i_24_1_48 XI2.XI1.XI14.XI3<7>.Y XI2.XI1.XI14.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<7>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<6>.MM_i_0 VSS! XI2.XI1.XI14.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<6>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<6>.MM_i_0_15 VSS! REG_DATA_2<6> XI2.XI1.XI14.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<6>.MM_i_0_15_63 XI2.XI1.XI14.XI3<6>.DUMMY1 REG_DATA_2<6>
+ XI2.XI1.XI14.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<6>.NEN
+ XI2.XI1.XI14.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<6>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<6>.MM_i_24 VDD! XI2.XI1.XI14.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<6>.MM_i_24_1 XI2.XI1.XI14.XI3<6>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<6>.MM_i_24_0 VDD! REG_DATA_2<6> XI2.XI1.XI14.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_2<6> XI2.XI1.XI14.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<6>.MM_i_24_1_48 XI2.XI1.XI14.XI3<6>.Y XI2.XI1.XI14.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<6>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<5>.MM_i_0 VSS! XI2.XI1.XI14.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<5>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<5>.MM_i_0_15 VSS! REG_DATA_2<5> XI2.XI1.XI14.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<5>.MM_i_0_15_63 XI2.XI1.XI14.XI3<5>.DUMMY1 REG_DATA_2<5>
+ XI2.XI1.XI14.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<5>.NEN
+ XI2.XI1.XI14.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<5>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<5>.MM_i_24 VDD! XI2.XI1.XI14.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<5>.MM_i_24_1 XI2.XI1.XI14.XI3<5>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<5>.MM_i_24_0 VDD! REG_DATA_2<5> XI2.XI1.XI14.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_2<5> XI2.XI1.XI14.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<5>.MM_i_24_1_48 XI2.XI1.XI14.XI3<5>.Y XI2.XI1.XI14.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<5>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<4>.MM_i_0 VSS! XI2.XI1.XI14.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<4>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<4>.MM_i_0_15 VSS! REG_DATA_2<4> XI2.XI1.XI14.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<4>.MM_i_0_15_63 XI2.XI1.XI14.XI3<4>.DUMMY1 REG_DATA_2<4>
+ XI2.XI1.XI14.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<4>.NEN
+ XI2.XI1.XI14.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<4>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<4>.MM_i_24 VDD! XI2.XI1.XI14.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<4>.MM_i_24_1 XI2.XI1.XI14.XI3<4>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<4>.MM_i_24_0 VDD! REG_DATA_2<4> XI2.XI1.XI14.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_2<4> XI2.XI1.XI14.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<4>.MM_i_24_1_48 XI2.XI1.XI14.XI3<4>.Y XI2.XI1.XI14.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<4>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<11>.MM_i_0 VSS! XI2.XI1.XI14.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<11>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<11>.MM_i_0_15 VSS! REG_DATA_2<11> XI2.XI1.XI14.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<11>.MM_i_0_15_63 XI2.XI1.XI14.XI3<11>.DUMMY1 REG_DATA_2<11>
+ XI2.XI1.XI14.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<11>.NEN
+ XI2.XI1.XI14.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<11>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<11>.MM_i_24 VDD! XI2.XI1.XI14.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<11>.MM_i_24_1 XI2.XI1.XI14.XI3<11>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<11>.MM_i_24_0 VDD! REG_DATA_2<11> XI2.XI1.XI14.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_2<11> XI2.XI1.XI14.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<11>.MM_i_24_1_48 XI2.XI1.XI14.XI3<11>.Y
+ XI2.XI1.XI14.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI14.XI3<11>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<10>.MM_i_0 VSS! XI2.XI1.XI14.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<10>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<10>.MM_i_0_15 VSS! REG_DATA_2<10> XI2.XI1.XI14.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<10>.MM_i_0_15_63 XI2.XI1.XI14.XI3<10>.DUMMY1 REG_DATA_2<10>
+ XI2.XI1.XI14.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<10>.NEN
+ XI2.XI1.XI14.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<10>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<10>.MM_i_24 VDD! XI2.XI1.XI14.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<10>.MM_i_24_1 XI2.XI1.XI14.XI3<10>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<10>.MM_i_24_0 VDD! REG_DATA_2<10> XI2.XI1.XI14.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_2<10> XI2.XI1.XI14.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<10>.MM_i_24_1_48 XI2.XI1.XI14.XI3<10>.Y
+ XI2.XI1.XI14.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI14.XI3<10>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<9>.MM_i_0 VSS! XI2.XI1.XI14.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<9>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<9>.MM_i_0_15 VSS! REG_DATA_2<9> XI2.XI1.XI14.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<9>.MM_i_0_15_63 XI2.XI1.XI14.XI3<9>.DUMMY1 REG_DATA_2<9>
+ XI2.XI1.XI14.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<9>.NEN
+ XI2.XI1.XI14.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<9>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<9>.MM_i_24 VDD! XI2.XI1.XI14.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<9>.MM_i_24_1 XI2.XI1.XI14.XI3<9>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<9>.MM_i_24_0 VDD! REG_DATA_2<9> XI2.XI1.XI14.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_2<9> XI2.XI1.XI14.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<9>.MM_i_24_1_48 XI2.XI1.XI14.XI3<9>.Y XI2.XI1.XI14.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<9>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<8>.MM_i_0 VSS! XI2.XI1.XI14.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<8>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<8>.MM_i_0_15 VSS! REG_DATA_2<8> XI2.XI1.XI14.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<8>.MM_i_0_15_63 XI2.XI1.XI14.XI3<8>.DUMMY1 REG_DATA_2<8>
+ XI2.XI1.XI14.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<8>.NEN
+ XI2.XI1.XI14.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<8>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<8>.MM_i_24 VDD! XI2.XI1.XI14.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<8>.MM_i_24_1 XI2.XI1.XI14.XI3<8>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<8>.MM_i_24_0 VDD! REG_DATA_2<8> XI2.XI1.XI14.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_2<8> XI2.XI1.XI14.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI14.XI3<8>.MM_i_24_1_48 XI2.XI1.XI14.XI3<8>.Y XI2.XI1.XI14.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI14.XI3<8>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<15>.MM_i_0 VSS! XI2.XI1.XI14.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<15>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<15>.MM_i_0_15 VSS! REG_DATA_2<15> XI2.XI1.XI14.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<15>.MM_i_0_15_63 XI2.XI1.XI14.XI3<15>.DUMMY1 REG_DATA_2<15>
+ XI2.XI1.XI14.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<15>.NEN
+ XI2.XI1.XI14.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<15>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<15>.MM_i_24 VDD! XI2.XI1.XI14.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<15>.MM_i_24_1 XI2.XI1.XI14.XI3<15>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<15>.MM_i_24_0 VDD! REG_DATA_2<15> XI2.XI1.XI14.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_2<15> XI2.XI1.XI14.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<15>.MM_i_24_1_48 XI2.XI1.XI14.XI3<15>.Y
+ XI2.XI1.XI14.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI14.XI3<15>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<14>.MM_i_0 VSS! XI2.XI1.XI14.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<14>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<14>.MM_i_0_15 VSS! REG_DATA_2<14> XI2.XI1.XI14.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<14>.MM_i_0_15_63 XI2.XI1.XI14.XI3<14>.DUMMY1 REG_DATA_2<14>
+ XI2.XI1.XI14.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<14>.NEN
+ XI2.XI1.XI14.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<14>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<14>.MM_i_24 VDD! XI2.XI1.XI14.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<14>.MM_i_24_1 XI2.XI1.XI14.XI3<14>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<14>.MM_i_24_0 VDD! REG_DATA_2<14> XI2.XI1.XI14.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_2<14> XI2.XI1.XI14.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<14>.MM_i_24_1_48 XI2.XI1.XI14.XI3<14>.Y
+ XI2.XI1.XI14.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI14.XI3<14>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<13>.MM_i_0 VSS! XI2.XI1.XI14.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<13>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<13>.MM_i_0_15 VSS! REG_DATA_2<13> XI2.XI1.XI14.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<13>.MM_i_0_15_63 XI2.XI1.XI14.XI3<13>.DUMMY1 REG_DATA_2<13>
+ XI2.XI1.XI14.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<13>.NEN
+ XI2.XI1.XI14.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<13>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<13>.MM_i_24 VDD! XI2.XI1.XI14.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<13>.MM_i_24_1 XI2.XI1.XI14.XI3<13>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<13>.MM_i_24_0 VDD! REG_DATA_2<13> XI2.XI1.XI14.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_2<13> XI2.XI1.XI14.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<13>.MM_i_24_1_48 XI2.XI1.XI14.XI3<13>.Y
+ XI2.XI1.XI14.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI14.XI3<13>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI14.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI14.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI14.XI3<12>.MM_i_0 VSS! XI2.XI1.XI14.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI14.XI3<12>.MM_i_0_14 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<12>.MM_i_0_15 VSS! REG_DATA_2<12> XI2.XI1.XI14.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<12>.MM_i_0_15_63 XI2.XI1.XI14.XI3<12>.DUMMY1 REG_DATA_2<12>
+ XI2.XI1.XI14.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI14.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI14.XI3<12>.NEN
+ XI2.XI1.XI14.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI14.XI3<12>.MM_i_17 VSS! XI2.NET1<10> XI2.XI1.XI14.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI14.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI14.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<12>.MM_i_24 VDD! XI2.XI1.XI14.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI14.XI3<12>.MM_i_24_1 XI2.XI1.XI14.XI3<12>.DUMMY0 XI2.NET1<10>
+ XI2.XI1.XI14.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI14.XI3<12>.MM_i_24_0 VDD! REG_DATA_2<12> XI2.XI1.XI14.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_2<12> XI2.XI1.XI14.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI14.XI3<12>.MM_i_24_1_48 XI2.XI1.XI14.XI3<12>.Y
+ XI2.XI1.XI14.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI14.XI3<12>.MM_i_42 VDD! XI2.NET1<10> XI2.XI1.XI14.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<3>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<3>.MM_i_0 VSS! XI2.XI1.XI13.XI3<3>.X RD_DATA_1<3> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<3>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<3>.MM_i_0_15 VSS! REG_DATA_1<3> XI2.XI1.XI13.XI3<3>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<3>.MM_i_0_15_63 XI2.XI1.XI13.XI3<3>.DUMMY1 REG_DATA_1<3>
+ XI2.XI1.XI13.XI3<3>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<3>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<3>.NEN
+ XI2.XI1.XI13.XI3<3>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<3>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<3>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<3>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<3>.MM_i_24 VDD! XI2.XI1.XI13.XI3<3>.Y RD_DATA_1<3> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<3>.MM_i_24_1 XI2.XI1.XI13.XI3<3>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<3>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<3>.MM_i_24_0 VDD! REG_DATA_1<3> XI2.XI1.XI13.XI3<3>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<3>.MM_i_24_0_64 VDD! REG_DATA_1<3> XI2.XI1.XI13.XI3<3>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<3>.MM_i_24_1_48 XI2.XI1.XI13.XI3<3>.Y XI2.XI1.XI13.XI3<3>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<3>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<3>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<2>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<2>.MM_i_0 VSS! XI2.XI1.XI13.XI3<2>.X RD_DATA_1<2> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<2>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<2>.MM_i_0_15 VSS! REG_DATA_1<2> XI2.XI1.XI13.XI3<2>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<2>.MM_i_0_15_63 XI2.XI1.XI13.XI3<2>.DUMMY1 REG_DATA_1<2>
+ XI2.XI1.XI13.XI3<2>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<2>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<2>.NEN
+ XI2.XI1.XI13.XI3<2>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<2>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<2>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<2>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<2>.MM_i_24 VDD! XI2.XI1.XI13.XI3<2>.Y RD_DATA_1<2> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<2>.MM_i_24_1 XI2.XI1.XI13.XI3<2>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<2>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<2>.MM_i_24_0 VDD! REG_DATA_1<2> XI2.XI1.XI13.XI3<2>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<2>.MM_i_24_0_64 VDD! REG_DATA_1<2> XI2.XI1.XI13.XI3<2>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<2>.MM_i_24_1_48 XI2.XI1.XI13.XI3<2>.Y XI2.XI1.XI13.XI3<2>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<2>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<2>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<1>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<1>.MM_i_0 VSS! XI2.XI1.XI13.XI3<1>.X RD_DATA_1<1> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<1>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<1>.MM_i_0_15 VSS! REG_DATA_1<1> XI2.XI1.XI13.XI3<1>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<1>.MM_i_0_15_63 XI2.XI1.XI13.XI3<1>.DUMMY1 REG_DATA_1<1>
+ XI2.XI1.XI13.XI3<1>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<1>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<1>.NEN
+ XI2.XI1.XI13.XI3<1>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<1>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<1>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<1>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<1>.MM_i_24 VDD! XI2.XI1.XI13.XI3<1>.Y RD_DATA_1<1> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<1>.MM_i_24_1 XI2.XI1.XI13.XI3<1>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<1>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<1>.MM_i_24_0 VDD! REG_DATA_1<1> XI2.XI1.XI13.XI3<1>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<1>.MM_i_24_0_64 VDD! REG_DATA_1<1> XI2.XI1.XI13.XI3<1>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<1>.MM_i_24_1_48 XI2.XI1.XI13.XI3<1>.Y XI2.XI1.XI13.XI3<1>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<1>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<1>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<0>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<0>.MM_i_0 VSS! XI2.XI1.XI13.XI3<0>.X RD_DATA_1<0> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<0>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<0>.MM_i_0_15 VSS! REG_DATA_1<0> XI2.XI1.XI13.XI3<0>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<0>.MM_i_0_15_63 XI2.XI1.XI13.XI3<0>.DUMMY1 REG_DATA_1<0>
+ XI2.XI1.XI13.XI3<0>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<0>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<0>.NEN
+ XI2.XI1.XI13.XI3<0>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<0>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<0>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<0>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<0>.MM_i_24 VDD! XI2.XI1.XI13.XI3<0>.Y RD_DATA_1<0> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<0>.MM_i_24_1 XI2.XI1.XI13.XI3<0>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<0>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<0>.MM_i_24_0 VDD! REG_DATA_1<0> XI2.XI1.XI13.XI3<0>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<0>.MM_i_24_0_64 VDD! REG_DATA_1<0> XI2.XI1.XI13.XI3<0>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<0>.MM_i_24_1_48 XI2.XI1.XI13.XI3<0>.Y XI2.XI1.XI13.XI3<0>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<0>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<0>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<7>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<7>.MM_i_0 VSS! XI2.XI1.XI13.XI3<7>.X RD_DATA_1<7> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<7>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<7>.MM_i_0_15 VSS! REG_DATA_1<7> XI2.XI1.XI13.XI3<7>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<7>.MM_i_0_15_63 XI2.XI1.XI13.XI3<7>.DUMMY1 REG_DATA_1<7>
+ XI2.XI1.XI13.XI3<7>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<7>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<7>.NEN
+ XI2.XI1.XI13.XI3<7>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<7>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<7>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<7>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<7>.MM_i_24 VDD! XI2.XI1.XI13.XI3<7>.Y RD_DATA_1<7> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<7>.MM_i_24_1 XI2.XI1.XI13.XI3<7>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<7>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<7>.MM_i_24_0 VDD! REG_DATA_1<7> XI2.XI1.XI13.XI3<7>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<7>.MM_i_24_0_64 VDD! REG_DATA_1<7> XI2.XI1.XI13.XI3<7>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<7>.MM_i_24_1_48 XI2.XI1.XI13.XI3<7>.Y XI2.XI1.XI13.XI3<7>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<7>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<7>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<6>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<6>.MM_i_0 VSS! XI2.XI1.XI13.XI3<6>.X RD_DATA_1<6> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<6>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<6>.MM_i_0_15 VSS! REG_DATA_1<6> XI2.XI1.XI13.XI3<6>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<6>.MM_i_0_15_63 XI2.XI1.XI13.XI3<6>.DUMMY1 REG_DATA_1<6>
+ XI2.XI1.XI13.XI3<6>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<6>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<6>.NEN
+ XI2.XI1.XI13.XI3<6>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<6>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<6>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<6>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<6>.MM_i_24 VDD! XI2.XI1.XI13.XI3<6>.Y RD_DATA_1<6> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<6>.MM_i_24_1 XI2.XI1.XI13.XI3<6>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<6>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<6>.MM_i_24_0 VDD! REG_DATA_1<6> XI2.XI1.XI13.XI3<6>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<6>.MM_i_24_0_64 VDD! REG_DATA_1<6> XI2.XI1.XI13.XI3<6>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<6>.MM_i_24_1_48 XI2.XI1.XI13.XI3<6>.Y XI2.XI1.XI13.XI3<6>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<6>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<6>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<5>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<5>.MM_i_0 VSS! XI2.XI1.XI13.XI3<5>.X RD_DATA_1<5> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<5>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<5>.MM_i_0_15 VSS! REG_DATA_1<5> XI2.XI1.XI13.XI3<5>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<5>.MM_i_0_15_63 XI2.XI1.XI13.XI3<5>.DUMMY1 REG_DATA_1<5>
+ XI2.XI1.XI13.XI3<5>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<5>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<5>.NEN
+ XI2.XI1.XI13.XI3<5>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<5>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<5>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<5>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<5>.MM_i_24 VDD! XI2.XI1.XI13.XI3<5>.Y RD_DATA_1<5> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<5>.MM_i_24_1 XI2.XI1.XI13.XI3<5>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<5>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<5>.MM_i_24_0 VDD! REG_DATA_1<5> XI2.XI1.XI13.XI3<5>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<5>.MM_i_24_0_64 VDD! REG_DATA_1<5> XI2.XI1.XI13.XI3<5>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<5>.MM_i_24_1_48 XI2.XI1.XI13.XI3<5>.Y XI2.XI1.XI13.XI3<5>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<5>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<5>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<4>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<4>.MM_i_0 VSS! XI2.XI1.XI13.XI3<4>.X RD_DATA_1<4> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<4>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<4>.MM_i_0_15 VSS! REG_DATA_1<4> XI2.XI1.XI13.XI3<4>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<4>.MM_i_0_15_63 XI2.XI1.XI13.XI3<4>.DUMMY1 REG_DATA_1<4>
+ XI2.XI1.XI13.XI3<4>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<4>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<4>.NEN
+ XI2.XI1.XI13.XI3<4>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<4>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<4>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<4>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<4>.MM_i_24 VDD! XI2.XI1.XI13.XI3<4>.Y RD_DATA_1<4> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<4>.MM_i_24_1 XI2.XI1.XI13.XI3<4>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<4>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<4>.MM_i_24_0 VDD! REG_DATA_1<4> XI2.XI1.XI13.XI3<4>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<4>.MM_i_24_0_64 VDD! REG_DATA_1<4> XI2.XI1.XI13.XI3<4>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<4>.MM_i_24_1_48 XI2.XI1.XI13.XI3<4>.Y XI2.XI1.XI13.XI3<4>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<4>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<4>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<11>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<11>.MM_i_0 VSS! XI2.XI1.XI13.XI3<11>.X RD_DATA_1<11> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<11>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<11>.MM_i_0_15 VSS! REG_DATA_1<11> XI2.XI1.XI13.XI3<11>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<11>.MM_i_0_15_63 XI2.XI1.XI13.XI3<11>.DUMMY1 REG_DATA_1<11>
+ XI2.XI1.XI13.XI3<11>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<11>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<11>.NEN
+ XI2.XI1.XI13.XI3<11>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<11>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<11>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<11>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<11>.MM_i_24 VDD! XI2.XI1.XI13.XI3<11>.Y RD_DATA_1<11> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<11>.MM_i_24_1 XI2.XI1.XI13.XI3<11>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<11>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<11>.MM_i_24_0 VDD! REG_DATA_1<11> XI2.XI1.XI13.XI3<11>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<11>.MM_i_24_0_64 VDD! REG_DATA_1<11> XI2.XI1.XI13.XI3<11>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<11>.MM_i_24_1_48 XI2.XI1.XI13.XI3<11>.Y
+ XI2.XI1.XI13.XI3<11>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI13.XI3<11>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<11>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<10>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<10>.MM_i_0 VSS! XI2.XI1.XI13.XI3<10>.X RD_DATA_1<10> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<10>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<10>.MM_i_0_15 VSS! REG_DATA_1<10> XI2.XI1.XI13.XI3<10>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<10>.MM_i_0_15_63 XI2.XI1.XI13.XI3<10>.DUMMY1 REG_DATA_1<10>
+ XI2.XI1.XI13.XI3<10>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<10>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<10>.NEN
+ XI2.XI1.XI13.XI3<10>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<10>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<10>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<10>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<10>.MM_i_24 VDD! XI2.XI1.XI13.XI3<10>.Y RD_DATA_1<10> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<10>.MM_i_24_1 XI2.XI1.XI13.XI3<10>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<10>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<10>.MM_i_24_0 VDD! REG_DATA_1<10> XI2.XI1.XI13.XI3<10>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<10>.MM_i_24_0_64 VDD! REG_DATA_1<10> XI2.XI1.XI13.XI3<10>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<10>.MM_i_24_1_48 XI2.XI1.XI13.XI3<10>.Y
+ XI2.XI1.XI13.XI3<10>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI13.XI3<10>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<10>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<9>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<9>.MM_i_0 VSS! XI2.XI1.XI13.XI3<9>.X RD_DATA_1<9> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<9>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<9>.MM_i_0_15 VSS! REG_DATA_1<9> XI2.XI1.XI13.XI3<9>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<9>.MM_i_0_15_63 XI2.XI1.XI13.XI3<9>.DUMMY1 REG_DATA_1<9>
+ XI2.XI1.XI13.XI3<9>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<9>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<9>.NEN
+ XI2.XI1.XI13.XI3<9>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<9>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<9>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<9>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<9>.MM_i_24 VDD! XI2.XI1.XI13.XI3<9>.Y RD_DATA_1<9> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<9>.MM_i_24_1 XI2.XI1.XI13.XI3<9>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<9>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<9>.MM_i_24_0 VDD! REG_DATA_1<9> XI2.XI1.XI13.XI3<9>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<9>.MM_i_24_0_64 VDD! REG_DATA_1<9> XI2.XI1.XI13.XI3<9>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<9>.MM_i_24_1_48 XI2.XI1.XI13.XI3<9>.Y XI2.XI1.XI13.XI3<9>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<9>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<9>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<8>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<8>.MM_i_0 VSS! XI2.XI1.XI13.XI3<8>.X RD_DATA_1<8> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<8>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<8>.MM_i_0_15 VSS! REG_DATA_1<8> XI2.XI1.XI13.XI3<8>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<8>.MM_i_0_15_63 XI2.XI1.XI13.XI3<8>.DUMMY1 REG_DATA_1<8>
+ XI2.XI1.XI13.XI3<8>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.22e-14
+ PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<8>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<8>.NEN
+ XI2.XI1.XI13.XI3<8>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<8>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<8>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<8>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<8>.MM_i_24 VDD! XI2.XI1.XI13.XI3<8>.Y RD_DATA_1<8> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<8>.MM_i_24_1 XI2.XI1.XI13.XI3<8>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<8>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14
+ PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<8>.MM_i_24_0 VDD! REG_DATA_1<8> XI2.XI1.XI13.XI3<8>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<8>.MM_i_24_0_64 VDD! REG_DATA_1<8> XI2.XI1.XI13.XI3<8>.Y VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI2.XI1.XI13.XI3<8>.MM_i_24_1_48 XI2.XI1.XI13.XI3<8>.Y XI2.XI1.XI13.XI3<8>.NEN
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06
+ PS=1.64e-06
mXI2.XI1.XI13.XI3<8>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<8>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<15>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<15>.MM_i_0 VSS! XI2.XI1.XI13.XI3<15>.X RD_DATA_1<15> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<15>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<15>.MM_i_0_15 VSS! REG_DATA_1<15> XI2.XI1.XI13.XI3<15>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<15>.MM_i_0_15_63 XI2.XI1.XI13.XI3<15>.DUMMY1 REG_DATA_1<15>
+ XI2.XI1.XI13.XI3<15>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<15>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<15>.NEN
+ XI2.XI1.XI13.XI3<15>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<15>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<15>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<15>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<15>.MM_i_24 VDD! XI2.XI1.XI13.XI3<15>.Y RD_DATA_1<15> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<15>.MM_i_24_1 XI2.XI1.XI13.XI3<15>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<15>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<15>.MM_i_24_0 VDD! REG_DATA_1<15> XI2.XI1.XI13.XI3<15>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<15>.MM_i_24_0_64 VDD! REG_DATA_1<15> XI2.XI1.XI13.XI3<15>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<15>.MM_i_24_1_48 XI2.XI1.XI13.XI3<15>.Y
+ XI2.XI1.XI13.XI3<15>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI13.XI3<15>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<15>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<14>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<14>.MM_i_0 VSS! XI2.XI1.XI13.XI3<14>.X RD_DATA_1<14> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<14>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<14>.MM_i_0_15 VSS! REG_DATA_1<14> XI2.XI1.XI13.XI3<14>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<14>.MM_i_0_15_63 XI2.XI1.XI13.XI3<14>.DUMMY1 REG_DATA_1<14>
+ XI2.XI1.XI13.XI3<14>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<14>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<14>.NEN
+ XI2.XI1.XI13.XI3<14>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<14>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<14>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<14>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<14>.MM_i_24 VDD! XI2.XI1.XI13.XI3<14>.Y RD_DATA_1<14> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<14>.MM_i_24_1 XI2.XI1.XI13.XI3<14>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<14>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<14>.MM_i_24_0 VDD! REG_DATA_1<14> XI2.XI1.XI13.XI3<14>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<14>.MM_i_24_0_64 VDD! REG_DATA_1<14> XI2.XI1.XI13.XI3<14>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<14>.MM_i_24_1_48 XI2.XI1.XI13.XI3<14>.Y
+ XI2.XI1.XI13.XI3<14>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI13.XI3<14>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<14>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<13>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<13>.MM_i_0 VSS! XI2.XI1.XI13.XI3<13>.X RD_DATA_1<13> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<13>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<13>.MM_i_0_15 VSS! REG_DATA_1<13> XI2.XI1.XI13.XI3<13>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<13>.MM_i_0_15_63 XI2.XI1.XI13.XI3<13>.DUMMY1 REG_DATA_1<13>
+ XI2.XI1.XI13.XI3<13>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<13>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<13>.NEN
+ XI2.XI1.XI13.XI3<13>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<13>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<13>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<13>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<13>.MM_i_24 VDD! XI2.XI1.XI13.XI3<13>.Y RD_DATA_1<13> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<13>.MM_i_24_1 XI2.XI1.XI13.XI3<13>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<13>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<13>.MM_i_24_0 VDD! REG_DATA_1<13> XI2.XI1.XI13.XI3<13>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<13>.MM_i_24_0_64 VDD! REG_DATA_1<13> XI2.XI1.XI13.XI3<13>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<13>.MM_i_24_1_48 XI2.XI1.XI13.XI3<13>.Y
+ XI2.XI1.XI13.XI3<13>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI13.XI3<13>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<13>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI2.XI1.XI13.XI3<12>.MM_i_0_6 VSS! XI2.XI1.XI13.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=3.7275e-14 AS=4.97e-14 PD=9.2e-07 PS=9.9e-07
mXI2.XI1.XI13.XI3<12>.MM_i_0 VSS! XI2.XI1.XI13.XI3<12>.X RD_DATA_1<12> VSS!
+ NMOS_VTL L=5e-08 W=3.55e-07 AD=9.4725e-14 AS=4.97e-14 PD=1.34e-06 PS=9.9e-07
mXI2.XI1.XI13.XI3<12>.MM_i_0_14 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=9.4725e-14 AS=5.81e-14 PD=1.34e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<12>.MM_i_0_15 VSS! REG_DATA_1<12> XI2.XI1.XI13.XI3<12>.X VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=3.22e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<12>.MM_i_0_15_63 XI2.XI1.XI13.XI3<12>.DUMMY1 REG_DATA_1<12>
+ XI2.XI1.XI13.XI3<12>.Y VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=3.22e-14 PD=1.11e-06 PS=1.04e-06
mXI2.XI1.XI13.XI3<12>.MM_i_0_14_47 VSS! XI2.XI1.XI13.XI3<12>.NEN
+ XI2.XI1.XI13.XI3<12>.DUMMY1 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI2.XI1.XI13.XI3<12>.MM_i_17 VSS! XI2.NET1<11> XI2.XI1.XI13.XI3<12>.NEN VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI2.XI1.XI13.XI3<12>.MM_i_24_3 VDD! XI2.XI1.XI13.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<12>.MM_i_24 VDD! XI2.XI1.XI13.XI3<12>.Y RD_DATA_1<12> VDD!
+ PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=7.56e-14 PD=1.29e-06 PS=1.36e-06
mXI2.XI1.XI13.XI3<12>.MM_i_24_1 XI2.XI1.XI13.XI3<12>.DUMMY0 XI2.NET1<11>
+ XI2.XI1.XI13.XI3<12>.X VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI2.XI1.XI13.XI3<12>.MM_i_24_0 VDD! REG_DATA_1<12> XI2.XI1.XI13.XI3<12>.DUMMY0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<12>.MM_i_24_0_64 VDD! REG_DATA_1<12> XI2.XI1.XI13.XI3<12>.Y
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI2.XI1.XI13.XI3<12>.MM_i_24_1_48 XI2.XI1.XI13.XI3<12>.Y
+ XI2.XI1.XI13.XI3<12>.NEN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.19e-14 PD=1.54e-06 PS=1.64e-06
mXI2.XI1.XI13.XI3<12>.MM_i_42 VDD! XI2.NET1<11> XI2.XI1.XI13.XI3<12>.NEN VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=3.3075e-14 PD=1.64e-06 PS=8.4e-07
mXI1.XI1.XI1.MM_i_0 XI1.XI1.WR_EN_BAR WR_EN VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI1.XI1.XI1.MM_i_1 XI1.XI1.WR_EN_BAR WR_EN VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI1.XI1.XI0.XI24.MM_i_1 XI1.XI1.XI0.XI24.NET_0 XI1.XI1.XI0.NET_11XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI24.MM_i_0 XI1.XI1.DEC_ADDR_BAR<12> XI1.XI1.XI0.NET_XX00
+ XI1.XI1.XI0.XI24.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI24.MM_i_3 XI1.XI1.DEC_ADDR_BAR<12> XI1.XI1.XI0.NET_11XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI24.MM_i_2 VDD! XI1.XI1.XI0.NET_XX00 XI1.XI1.DEC_ADDR_BAR<12> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI23.MM_i_1 XI1.XI1.XI0.XI23.NET_0 XI1.XI1.XI0.NET_10XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI23.MM_i_0 XI1.XI1.DEC_ADDR_BAR<11> XI1.XI1.XI0.NET_XX11
+ XI1.XI1.XI0.XI23.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI23.MM_i_3 XI1.XI1.DEC_ADDR_BAR<11> XI1.XI1.XI0.NET_10XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI23.MM_i_2 VDD! XI1.XI1.XI0.NET_XX11 XI1.XI1.DEC_ADDR_BAR<11> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI22.MM_i_1 XI1.XI1.XI0.XI22.NET_0 XI1.XI1.XI0.NET_10XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI22.MM_i_0 XI1.XI1.DEC_ADDR_BAR<10> XI1.XI1.XI0.NET_XX10
+ XI1.XI1.XI0.XI22.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI22.MM_i_3 XI1.XI1.DEC_ADDR_BAR<10> XI1.XI1.XI0.NET_10XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI22.MM_i_2 VDD! XI1.XI1.XI0.NET_XX10 XI1.XI1.DEC_ADDR_BAR<10> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI21.MM_i_1 XI1.XI1.XI0.XI21.NET_0 XI1.XI1.XI0.NET_10XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI21.MM_i_0 XI1.XI1.DEC_ADDR_BAR<9> XI1.XI1.XI0.NET_XX01
+ XI1.XI1.XI0.XI21.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI21.MM_i_3 XI1.XI1.DEC_ADDR_BAR<9> XI1.XI1.XI0.NET_10XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI21.MM_i_2 VDD! XI1.XI1.XI0.NET_XX01 XI1.XI1.DEC_ADDR_BAR<9> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI20.MM_i_1 XI1.XI1.XI0.XI20.NET_0 XI1.XI1.XI0.NET_10XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI20.MM_i_0 XI1.XI1.DEC_ADDR_BAR<8> XI1.XI1.XI0.NET_XX00
+ XI1.XI1.XI0.XI20.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI20.MM_i_3 XI1.XI1.DEC_ADDR_BAR<8> XI1.XI1.XI0.NET_10XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI20.MM_i_2 VDD! XI1.XI1.XI0.NET_XX00 XI1.XI1.DEC_ADDR_BAR<8> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI19.MM_i_1 XI1.XI1.XI0.XI19.NET_0 XI1.XI1.XI0.NET_01XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI19.MM_i_0 XI1.XI1.DEC_ADDR_BAR<7> XI1.XI1.XI0.NET_XX11
+ XI1.XI1.XI0.XI19.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI19.MM_i_3 XI1.XI1.DEC_ADDR_BAR<7> XI1.XI1.XI0.NET_01XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI19.MM_i_2 VDD! XI1.XI1.XI0.NET_XX11 XI1.XI1.DEC_ADDR_BAR<7> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI18.MM_i_1 XI1.XI1.XI0.XI18.NET_0 XI1.XI1.XI0.NET_01XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI18.MM_i_0 XI1.XI1.DEC_ADDR_BAR<6> XI1.XI1.XI0.NET_XX10
+ XI1.XI1.XI0.XI18.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI18.MM_i_3 XI1.XI1.DEC_ADDR_BAR<6> XI1.XI1.XI0.NET_01XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI18.MM_i_2 VDD! XI1.XI1.XI0.NET_XX10 XI1.XI1.DEC_ADDR_BAR<6> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI17.MM_i_1 XI1.XI1.XI0.XI17.NET_0 XI1.XI1.XI0.NET_01XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI17.MM_i_0 XI1.XI1.DEC_ADDR_BAR<5> XI1.XI1.XI0.NET_XX01
+ XI1.XI1.XI0.XI17.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI17.MM_i_3 XI1.XI1.DEC_ADDR_BAR<5> XI1.XI1.XI0.NET_01XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI17.MM_i_2 VDD! XI1.XI1.XI0.NET_XX01 XI1.XI1.DEC_ADDR_BAR<5> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI16.MM_i_1 XI1.XI1.XI0.XI16.NET_0 XI1.XI1.XI0.NET_01XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI16.MM_i_0 XI1.XI1.DEC_ADDR_BAR<4> XI1.XI1.XI0.NET_XX00
+ XI1.XI1.XI0.XI16.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI16.MM_i_3 XI1.XI1.DEC_ADDR_BAR<4> XI1.XI1.XI0.NET_01XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI16.MM_i_2 VDD! XI1.XI1.XI0.NET_XX00 XI1.XI1.DEC_ADDR_BAR<4> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI15.MM_i_1 XI1.XI1.XI0.XI15.NET_0 XI1.XI1.XI0.NET_00XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI15.MM_i_0 XI1.XI1.DEC_ADDR_BAR<3> XI1.XI1.XI0.NET_XX11
+ XI1.XI1.XI0.XI15.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI15.MM_i_3 XI1.XI1.DEC_ADDR_BAR<3> XI1.XI1.XI0.NET_00XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI15.MM_i_2 VDD! XI1.XI1.XI0.NET_XX11 XI1.XI1.DEC_ADDR_BAR<3> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI14.MM_i_1 XI1.XI1.XI0.XI14.NET_0 XI1.XI1.XI0.NET_00XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI14.MM_i_0 XI1.XI1.DEC_ADDR_BAR<2> XI1.XI1.XI0.NET_XX10
+ XI1.XI1.XI0.XI14.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI14.MM_i_3 XI1.XI1.DEC_ADDR_BAR<2> XI1.XI1.XI0.NET_00XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI14.MM_i_2 VDD! XI1.XI1.XI0.NET_XX10 XI1.XI1.DEC_ADDR_BAR<2> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI13.MM_i_1 XI1.XI1.XI0.XI13.NET_0 XI1.XI1.XI0.NET_00XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI13.MM_i_0 XI1.XI1.DEC_ADDR_BAR<1> XI1.XI1.XI0.NET_XX01
+ XI1.XI1.XI0.XI13.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI13.MM_i_3 XI1.XI1.DEC_ADDR_BAR<1> XI1.XI1.XI0.NET_00XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI13.MM_i_2 VDD! XI1.XI1.XI0.NET_XX01 XI1.XI1.DEC_ADDR_BAR<1> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI12.MM_i_1 XI1.XI1.XI0.XI12.NET_0 XI1.XI1.XI0.NET_00XX VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI0.XI12.MM_i_0 XI1.XI1.DEC_ADDR_BAR<0> XI1.XI1.XI0.NET_XX00
+ XI1.XI1.XI0.XI12.NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI12.MM_i_3 XI1.XI1.DEC_ADDR_BAR<0> XI1.XI1.XI0.NET_00XX VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI0.XI12.MM_i_2 VDD! XI1.XI1.XI0.NET_XX00 XI1.XI1.DEC_ADDR_BAR<0> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI11.MM_i_2 XI1.XI1.XI0.XI11.NET_0 WR_ADDR<2>
+ XI1.XI1.XI0.XI11.ZN_NEG VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI11.MM_i_3 VSS! WR_ADDR<3> XI1.XI1.XI0.XI11.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI11.MM_i_0 XI1.XI1.XI0.NET_11XX XI1.XI1.XI0.XI11.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI11.MM_i_4 XI1.XI1.XI0.XI11.ZN_NEG WR_ADDR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI11.MM_i_5 VDD! WR_ADDR<3> XI1.XI1.XI0.XI11.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI11.MM_i_1 XI1.XI1.XI0.NET_11XX XI1.XI1.XI0.XI11.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI7.MM_i_2 XI1.XI1.XI0.XI7.NET_0 WR_ADDR<0> XI1.XI1.XI0.XI7.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI7.MM_i_3 VSS! WR_ADDR<1> XI1.XI1.XI0.XI7.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI7.MM_i_0 XI1.XI1.XI0.NET_XX11 XI1.XI1.XI0.XI7.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI7.MM_i_4 XI1.XI1.XI0.XI7.ZN_NEG WR_ADDR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI7.MM_i_5 VDD! WR_ADDR<1> XI1.XI1.XI0.XI7.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI7.MM_i_1 XI1.XI1.XI0.NET_XX11 XI1.XI1.XI0.XI7.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI10.MM_i_2 XI1.XI1.XI0.XI10.NET_0 XI1.XI1.XI0.ADDR_BAR<2>
+ XI1.XI1.XI0.XI10.ZN_NEG VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI10.MM_i_3 VSS! WR_ADDR<3> XI1.XI1.XI0.XI10.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI10.MM_i_0 XI1.XI1.XI0.NET_10XX XI1.XI1.XI0.XI10.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI10.MM_i_4 XI1.XI1.XI0.XI10.ZN_NEG XI1.XI1.XI0.ADDR_BAR<2> VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI1.XI0.XI10.MM_i_5 VDD! WR_ADDR<3> XI1.XI1.XI0.XI10.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI10.MM_i_1 XI1.XI1.XI0.NET_10XX XI1.XI1.XI0.XI10.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI6.MM_i_2 XI1.XI1.XI0.XI6.NET_0 XI1.XI1.XI0.ADDR_BAR<0>
+ XI1.XI1.XI0.XI6.ZN_NEG VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI6.MM_i_3 VSS! WR_ADDR<1> XI1.XI1.XI0.XI6.NET_0 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI6.MM_i_0 XI1.XI1.XI0.NET_XX10 XI1.XI1.XI0.XI6.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI6.MM_i_4 XI1.XI1.XI0.XI6.ZN_NEG XI1.XI1.XI0.ADDR_BAR<0> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI6.MM_i_5 VDD! WR_ADDR<1> XI1.XI1.XI0.XI6.ZN_NEG VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI6.MM_i_1 XI1.XI1.XI0.NET_XX10 XI1.XI1.XI0.XI6.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI9.MM_i_2 XI1.XI1.XI0.XI9.NET_0 WR_ADDR<2> XI1.XI1.XI0.XI9.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI9.MM_i_3 VSS! XI1.XI1.XI0.ADDR_BAR<3> XI1.XI1.XI0.XI9.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI9.MM_i_0 XI1.XI1.XI0.NET_01XX XI1.XI1.XI0.XI9.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI9.MM_i_4 XI1.XI1.XI0.XI9.ZN_NEG WR_ADDR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI9.MM_i_5 VDD! XI1.XI1.XI0.ADDR_BAR<3> XI1.XI1.XI0.XI9.ZN_NEG VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI9.MM_i_1 XI1.XI1.XI0.NET_01XX XI1.XI1.XI0.XI9.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI5.MM_i_2 XI1.XI1.XI0.XI5.NET_0 WR_ADDR<0> XI1.XI1.XI0.XI5.ZN_NEG
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI5.MM_i_3 VSS! XI1.XI1.XI0.ADDR_BAR<1> XI1.XI1.XI0.XI5.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI5.MM_i_0 XI1.XI1.XI0.NET_XX01 XI1.XI1.XI0.XI5.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI5.MM_i_4 XI1.XI1.XI0.XI5.ZN_NEG WR_ADDR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI5.MM_i_5 VDD! XI1.XI1.XI0.ADDR_BAR<1> XI1.XI1.XI0.XI5.ZN_NEG VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI5.MM_i_1 XI1.XI1.XI0.NET_XX01 XI1.XI1.XI0.XI5.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI8.MM_i_2 XI1.XI1.XI0.XI8.NET_0 XI1.XI1.XI0.ADDR_BAR<2>
+ XI1.XI1.XI0.XI8.ZN_NEG VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI8.MM_i_3 VSS! XI1.XI1.XI0.ADDR_BAR<3> XI1.XI1.XI0.XI8.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI8.MM_i_0 XI1.XI1.XI0.NET_00XX XI1.XI1.XI0.XI8.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI8.MM_i_4 XI1.XI1.XI0.XI8.ZN_NEG XI1.XI1.XI0.ADDR_BAR<2> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI8.MM_i_5 VDD! XI1.XI1.XI0.ADDR_BAR<3> XI1.XI1.XI0.XI8.ZN_NEG VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI8.MM_i_1 XI1.XI1.XI0.NET_00XX XI1.XI1.XI0.XI8.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI4.MM_i_2 XI1.XI1.XI0.XI4.NET_0 XI1.XI1.XI0.ADDR_BAR<0>
+ XI1.XI1.XI0.XI4.ZN_NEG VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI1.XI0.XI4.MM_i_3 VSS! XI1.XI1.XI0.ADDR_BAR<1> XI1.XI1.XI0.XI4.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI1.XI1.XI0.XI4.MM_i_0 XI1.XI1.XI0.NET_XX00 XI1.XI1.XI0.XI4.ZN_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI0.XI4.MM_i_4 XI1.XI1.XI0.XI4.ZN_NEG XI1.XI1.XI0.ADDR_BAR<0> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI1.XI0.XI4.MM_i_5 VDD! XI1.XI1.XI0.ADDR_BAR<1> XI1.XI1.XI0.XI4.ZN_NEG VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI1.XI1.XI0.XI4.MM_i_1 XI1.XI1.XI0.NET_XX00 XI1.XI1.XI0.XI4.ZN_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI0.XI2.MM_i_0 XI1.XI1.XI0.ADDR_BAR<2> WR_ADDR<2> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI1.XI1.XI0.XI2.MM_i_1 XI1.XI1.XI0.ADDR_BAR<2> WR_ADDR<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI1.XI1.XI0.XI0.MM_i_0 XI1.XI1.XI0.ADDR_BAR<0> WR_ADDR<0> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI1.XI1.XI0.XI0.MM_i_1 XI1.XI1.XI0.ADDR_BAR<0> WR_ADDR<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI1.XI1.XI0.XI3.MM_i_0 XI1.XI1.XI0.ADDR_BAR<3> WR_ADDR<3> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI1.XI1.XI0.XI3.MM_i_1 XI1.XI1.XI0.ADDR_BAR<3> WR_ADDR<3> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI1.XI1.XI0.XI1.MM_i_0 XI1.XI1.XI0.ADDR_BAR<1> WR_ADDR<1> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI1.XI1.XI0.XI1.MM_i_1 XI1.XI1.XI0.ADDR_BAR<1> WR_ADDR<1> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI1.XI1.XI2<12>.MM_i_1 XI1.WR_ADDR_EN<12> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<12>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<12> XI1.WR_ADDR_EN<12> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<12>.MM_i_3 XI1.XI1.XI2<12>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<12>.MM_i_2 XI1.WR_ADDR_EN<12> XI1.XI1.DEC_ADDR_BAR<12>
+ XI1.XI1.XI2<12>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<11>.MM_i_1 XI1.WR_ADDR_EN<11> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<11>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<11> XI1.WR_ADDR_EN<11> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<11>.MM_i_3 XI1.XI1.XI2<11>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<11>.MM_i_2 XI1.WR_ADDR_EN<11> XI1.XI1.DEC_ADDR_BAR<11>
+ XI1.XI1.XI2<11>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<10>.MM_i_1 XI1.WR_ADDR_EN<10> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<10>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<10> XI1.WR_ADDR_EN<10> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<10>.MM_i_3 XI1.XI1.XI2<10>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<10>.MM_i_2 XI1.WR_ADDR_EN<10> XI1.XI1.DEC_ADDR_BAR<10>
+ XI1.XI1.XI2<10>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<9>.MM_i_1 XI1.WR_ADDR_EN<9> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<9>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<9> XI1.WR_ADDR_EN<9> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<9>.MM_i_3 XI1.XI1.XI2<9>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<9>.MM_i_2 XI1.WR_ADDR_EN<9> XI1.XI1.DEC_ADDR_BAR<9>
+ XI1.XI1.XI2<9>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<8>.MM_i_1 XI1.WR_ADDR_EN<8> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<8>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<8> XI1.WR_ADDR_EN<8> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<8>.MM_i_3 XI1.XI1.XI2<8>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<8>.MM_i_2 XI1.WR_ADDR_EN<8> XI1.XI1.DEC_ADDR_BAR<8>
+ XI1.XI1.XI2<8>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<7>.MM_i_1 XI1.WR_ADDR_EN<7> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<7>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<7> XI1.WR_ADDR_EN<7> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<7>.MM_i_3 XI1.XI1.XI2<7>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<7>.MM_i_2 XI1.WR_ADDR_EN<7> XI1.XI1.DEC_ADDR_BAR<7>
+ XI1.XI1.XI2<7>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<6>.MM_i_1 XI1.WR_ADDR_EN<6> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<6>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<6> XI1.WR_ADDR_EN<6> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<6>.MM_i_3 XI1.XI1.XI2<6>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<6>.MM_i_2 XI1.WR_ADDR_EN<6> XI1.XI1.DEC_ADDR_BAR<6>
+ XI1.XI1.XI2<6>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<5>.MM_i_1 XI1.WR_ADDR_EN<5> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<5>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<5> XI1.WR_ADDR_EN<5> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<5>.MM_i_3 XI1.XI1.XI2<5>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<5>.MM_i_2 XI1.WR_ADDR_EN<5> XI1.XI1.DEC_ADDR_BAR<5>
+ XI1.XI1.XI2<5>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<4>.MM_i_1 XI1.WR_ADDR_EN<4> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<4>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<4> XI1.WR_ADDR_EN<4> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<4>.MM_i_3 XI1.XI1.XI2<4>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<4>.MM_i_2 XI1.WR_ADDR_EN<4> XI1.XI1.DEC_ADDR_BAR<4>
+ XI1.XI1.XI2<4>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<3>.MM_i_1 XI1.WR_ADDR_EN<3> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<3>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<3> XI1.WR_ADDR_EN<3> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<3>.MM_i_3 XI1.XI1.XI2<3>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<3>.MM_i_2 XI1.WR_ADDR_EN<3> XI1.XI1.DEC_ADDR_BAR<3>
+ XI1.XI1.XI2<3>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<2>.MM_i_1 XI1.WR_ADDR_EN<2> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<2>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<2> XI1.WR_ADDR_EN<2> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<2>.MM_i_3 XI1.XI1.XI2<2>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<2>.MM_i_2 XI1.WR_ADDR_EN<2> XI1.XI1.DEC_ADDR_BAR<2>
+ XI1.XI1.XI2<2>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<1>.MM_i_1 XI1.WR_ADDR_EN<1> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<1>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<1> XI1.WR_ADDR_EN<1> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<1>.MM_i_3 XI1.XI1.XI2<1>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<1>.MM_i_2 XI1.WR_ADDR_EN<1> XI1.XI1.DEC_ADDR_BAR<1>
+ XI1.XI1.XI2<1>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI1.XI2<0>.MM_i_1 XI1.WR_ADDR_EN<0> XI1.XI1.WR_EN_BAR VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI1.XI2<0>.MM_i_0 VSS! XI1.XI1.DEC_ADDR_BAR<0> XI1.WR_ADDR_EN<0> VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI1.XI2<0>.MM_i_3 XI1.XI1.XI2<0>.NET_0 XI1.XI1.WR_EN_BAR VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI1.XI2<0>.MM_i_2 XI1.WR_ADDR_EN<0> XI1.XI1.DEC_ADDR_BAR<0>
+ XI1.XI1.XI2<0>.NET_0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14
+ PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI18.MM_i_0 VSS! XI1.XI0.CK_EN<3> XI1.XI0.NET18 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI18.MM_i_1 XI1.XI0.NET18 XI1.XI0.CK_EN<2> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI18.MM_i_2 VSS! XI1.XI0.CK_EN<1> XI1.XI0.NET18 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI18.MM_i_3 XI1.XI0.NET18 XI1.XI0.CK_EN<0> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI19.MM_i_0 XI1.XI0.CLK_PREBUFF XI1.XI0.NET9 XI1.XI0.XI19.NET_0 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI19.MM_i_1 XI1.XI0.XI19.NET_0 XI1.XI0.NET5 XI1.XI0.XI19.NET_1 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI19.MM_i_2 XI1.XI0.XI19.NET_1 XI1.XI0.NET13 XI1.XI0.XI19.NET_2 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI19.MM_i_3 XI1.XI0.XI19.NET_2 XI1.XI0.NET18 VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI18.MM_i_4 XI1.XI0.NET18 XI1.XI0.CK_EN<3> XI1.XI0.XI18.NET_0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI18.MM_i_5 XI1.XI0.XI18.NET_0 XI1.XI0.CK_EN<2> XI1.XI0.XI18.NET_1 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI18.MM_i_6 XI1.XI0.XI18.NET_1 XI1.XI0.CK_EN<1> XI1.XI0.XI18.NET_2 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI18.MM_i_7 XI1.XI0.XI18.NET_2 XI1.XI0.CK_EN<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI19.MM_i_4 VDD! XI1.XI0.NET9 XI1.XI0.CLK_PREBUFF VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI19.MM_i_5 XI1.XI0.CLK_PREBUFF XI1.XI0.NET5 VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI19.MM_i_6 VDD! XI1.XI0.NET13 XI1.XI0.CLK_PREBUFF VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI19.MM_i_7 XI1.XI0.CLK_PREBUFF XI1.XI0.NET18 VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<12>.MM_i_0 VSS! XI1.XI0.XI14<12>.NET_002 XI1.XI0.XI14<12>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<12>.MM_i_21 VSS! XI1.WR_ADDR_EN<12> XI1.XI0.XI14<12>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<12>.MM_i_17 XI1.XI0.XI14<12>.NET_003 XI1.XI0.XI14<12>.NET_005
+ XI1.XI0.XI14<12>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<12>.MM_i_11 XI1.XI0.XI14<12>.NET_002 XI1.XI0.XI14<12>.NET_004
+ XI1.XI0.XI14<12>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<12>.MM_i_7 XI1.XI0.XI14<12>.NET_001 XI1.XI0.XI14<12>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<12>.MM_i_27 XI1.XI0.XI14<12>.NET_004 XI1.XI0.XI14<12>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<12>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<12>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<12>.MM_i_40 XI1.XI0.XI14<12>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<12>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<12>.MM_i_45 VSS! XI1.XI0.XI14<12>.NET_000 XI1.XI0.XI14<12>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<12>.MM_i_51 XI1.XI0.CK_EN<12> XI1.XI0.XI14<12>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<12>.MM_i_51_7 XI1.XI0.CK_EN<12> XI1.XI0.XI14<12>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<12>.MM_i_57 VDD! XI1.XI0.XI14<12>.NET_002 XI1.XI0.XI14<12>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<12>.MM_i_78 VDD! XI1.WR_ADDR_EN<12> XI1.XI0.XI14<12>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<12>.MM_i_74 XI1.XI0.XI14<12>.NET_009 XI1.XI0.XI14<12>.NET_004
+ XI1.XI0.XI14<12>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<12>.MM_i_68 XI1.XI0.XI14<12>.NET_002 XI1.XI0.XI14<12>.NET_005
+ XI1.XI0.XI14<12>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<12>.MM_i_64 XI1.XI0.XI14<12>.NET_008 XI1.XI0.XI14<12>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<12>.MM_i_84 XI1.XI0.XI14<12>.NET_004 XI1.XI0.XI14<12>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<12>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<12>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<12>.MM_i_97 XI1.XI0.XI14<12>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<12>.MM_i_103 VDD! XI1.XI0.XI14<12>.NET_000
+ XI1.XI0.XI14<12>.NET_006 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13
+ AS=8.82e-14 PD=1.59e-06 PS=1.54e-06
mXI1.XI0.XI14<12>.MM_i_109 XI1.XI0.CK_EN<12> XI1.XI0.XI14<12>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<12>.MM_i_109_4 XI1.XI0.CK_EN<12> XI1.XI0.XI14<12>.NET_006 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06
+ PS=1.47e-06
mXI1.XI0.XI14<11>.MM_i_0 VSS! XI1.XI0.XI14<11>.NET_002 XI1.XI0.XI14<11>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<11>.MM_i_21 VSS! XI1.WR_ADDR_EN<11> XI1.XI0.XI14<11>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<11>.MM_i_17 XI1.XI0.XI14<11>.NET_003 XI1.XI0.XI14<11>.NET_005
+ XI1.XI0.XI14<11>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<11>.MM_i_11 XI1.XI0.XI14<11>.NET_002 XI1.XI0.XI14<11>.NET_004
+ XI1.XI0.XI14<11>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<11>.MM_i_7 XI1.XI0.XI14<11>.NET_001 XI1.XI0.XI14<11>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<11>.MM_i_27 XI1.XI0.XI14<11>.NET_004 XI1.XI0.XI14<11>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<11>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<11>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<11>.MM_i_40 XI1.XI0.XI14<11>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<11>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<11>.MM_i_45 VSS! XI1.XI0.XI14<11>.NET_000 XI1.XI0.XI14<11>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<11>.MM_i_51 XI1.XI0.CK_EN<11> XI1.XI0.XI14<11>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<11>.MM_i_51_7 XI1.XI0.CK_EN<11> XI1.XI0.XI14<11>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<11>.MM_i_57 VDD! XI1.XI0.XI14<11>.NET_002 XI1.XI0.XI14<11>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<11>.MM_i_78 VDD! XI1.WR_ADDR_EN<11> XI1.XI0.XI14<11>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<11>.MM_i_74 XI1.XI0.XI14<11>.NET_009 XI1.XI0.XI14<11>.NET_004
+ XI1.XI0.XI14<11>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<11>.MM_i_68 XI1.XI0.XI14<11>.NET_002 XI1.XI0.XI14<11>.NET_005
+ XI1.XI0.XI14<11>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<11>.MM_i_64 XI1.XI0.XI14<11>.NET_008 XI1.XI0.XI14<11>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<11>.MM_i_84 XI1.XI0.XI14<11>.NET_004 XI1.XI0.XI14<11>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<11>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<11>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<11>.MM_i_97 XI1.XI0.XI14<11>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<11>.MM_i_103 VDD! XI1.XI0.XI14<11>.NET_000
+ XI1.XI0.XI14<11>.NET_006 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13
+ AS=8.82e-14 PD=1.59e-06 PS=1.54e-06
mXI1.XI0.XI14<11>.MM_i_109 XI1.XI0.CK_EN<11> XI1.XI0.XI14<11>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<11>.MM_i_109_4 XI1.XI0.CK_EN<11> XI1.XI0.XI14<11>.NET_006 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06
+ PS=1.47e-06
mXI1.XI0.XI14<10>.MM_i_0 VSS! XI1.XI0.XI14<10>.NET_002 XI1.XI0.XI14<10>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<10>.MM_i_21 VSS! XI1.WR_ADDR_EN<10> XI1.XI0.XI14<10>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<10>.MM_i_17 XI1.XI0.XI14<10>.NET_003 XI1.XI0.XI14<10>.NET_005
+ XI1.XI0.XI14<10>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<10>.MM_i_11 XI1.XI0.XI14<10>.NET_002 XI1.XI0.XI14<10>.NET_004
+ XI1.XI0.XI14<10>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<10>.MM_i_7 XI1.XI0.XI14<10>.NET_001 XI1.XI0.XI14<10>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<10>.MM_i_27 XI1.XI0.XI14<10>.NET_004 XI1.XI0.XI14<10>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<10>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<10>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<10>.MM_i_40 XI1.XI0.XI14<10>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<10>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<10>.MM_i_45 VSS! XI1.XI0.XI14<10>.NET_000 XI1.XI0.XI14<10>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<10>.MM_i_51 XI1.XI0.CK_EN<10> XI1.XI0.XI14<10>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<10>.MM_i_51_7 XI1.XI0.CK_EN<10> XI1.XI0.XI14<10>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<10>.MM_i_57 VDD! XI1.XI0.XI14<10>.NET_002 XI1.XI0.XI14<10>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<10>.MM_i_78 VDD! XI1.WR_ADDR_EN<10> XI1.XI0.XI14<10>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<10>.MM_i_74 XI1.XI0.XI14<10>.NET_009 XI1.XI0.XI14<10>.NET_004
+ XI1.XI0.XI14<10>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<10>.MM_i_68 XI1.XI0.XI14<10>.NET_002 XI1.XI0.XI14<10>.NET_005
+ XI1.XI0.XI14<10>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<10>.MM_i_64 XI1.XI0.XI14<10>.NET_008 XI1.XI0.XI14<10>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<10>.MM_i_84 XI1.XI0.XI14<10>.NET_004 XI1.XI0.XI14<10>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<10>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<10>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<10>.MM_i_97 XI1.XI0.XI14<10>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<10>.MM_i_103 VDD! XI1.XI0.XI14<10>.NET_000
+ XI1.XI0.XI14<10>.NET_006 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13
+ AS=8.82e-14 PD=1.59e-06 PS=1.54e-06
mXI1.XI0.XI14<10>.MM_i_109 XI1.XI0.CK_EN<10> XI1.XI0.XI14<10>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<10>.MM_i_109_4 XI1.XI0.CK_EN<10> XI1.XI0.XI14<10>.NET_006 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06
+ PS=1.47e-06
mXI1.XI0.XI14<9>.MM_i_0 VSS! XI1.XI0.XI14<9>.NET_002 XI1.XI0.XI14<9>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<9>.MM_i_21 VSS! XI1.WR_ADDR_EN<9> XI1.XI0.XI14<9>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<9>.MM_i_17 XI1.XI0.XI14<9>.NET_003 XI1.XI0.XI14<9>.NET_005
+ XI1.XI0.XI14<9>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<9>.MM_i_11 XI1.XI0.XI14<9>.NET_002 XI1.XI0.XI14<9>.NET_004
+ XI1.XI0.XI14<9>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<9>.MM_i_7 XI1.XI0.XI14<9>.NET_001 XI1.XI0.XI14<9>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<9>.MM_i_27 XI1.XI0.XI14<9>.NET_004 XI1.XI0.XI14<9>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<9>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<9>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<9>.MM_i_40 XI1.XI0.XI14<9>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<9>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<9>.MM_i_45 VSS! XI1.XI0.XI14<9>.NET_000 XI1.XI0.XI14<9>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<9>.MM_i_51 XI1.XI0.CK_EN<9> XI1.XI0.XI14<9>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<9>.MM_i_51_7 XI1.XI0.CK_EN<9> XI1.XI0.XI14<9>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<9>.MM_i_57 VDD! XI1.XI0.XI14<9>.NET_002 XI1.XI0.XI14<9>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<9>.MM_i_78 VDD! XI1.WR_ADDR_EN<9> XI1.XI0.XI14<9>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<9>.MM_i_74 XI1.XI0.XI14<9>.NET_009 XI1.XI0.XI14<9>.NET_004
+ XI1.XI0.XI14<9>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<9>.MM_i_68 XI1.XI0.XI14<9>.NET_002 XI1.XI0.XI14<9>.NET_005
+ XI1.XI0.XI14<9>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<9>.MM_i_64 XI1.XI0.XI14<9>.NET_008 XI1.XI0.XI14<9>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<9>.MM_i_84 XI1.XI0.XI14<9>.NET_004 XI1.XI0.XI14<9>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<9>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<9>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<9>.MM_i_97 XI1.XI0.XI14<9>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<9>.MM_i_103 VDD! XI1.XI0.XI14<9>.NET_000 XI1.XI0.XI14<9>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<9>.MM_i_109 XI1.XI0.CK_EN<9> XI1.XI0.XI14<9>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<9>.MM_i_109_4 XI1.XI0.CK_EN<9> XI1.XI0.XI14<9>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<8>.MM_i_0 VSS! XI1.XI0.XI14<8>.NET_002 XI1.XI0.XI14<8>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<8>.MM_i_21 VSS! XI1.WR_ADDR_EN<8> XI1.XI0.XI14<8>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<8>.MM_i_17 XI1.XI0.XI14<8>.NET_003 XI1.XI0.XI14<8>.NET_005
+ XI1.XI0.XI14<8>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<8>.MM_i_11 XI1.XI0.XI14<8>.NET_002 XI1.XI0.XI14<8>.NET_004
+ XI1.XI0.XI14<8>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<8>.MM_i_7 XI1.XI0.XI14<8>.NET_001 XI1.XI0.XI14<8>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<8>.MM_i_27 XI1.XI0.XI14<8>.NET_004 XI1.XI0.XI14<8>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<8>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<8>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<8>.MM_i_40 XI1.XI0.XI14<8>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<8>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<8>.MM_i_45 VSS! XI1.XI0.XI14<8>.NET_000 XI1.XI0.XI14<8>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<8>.MM_i_51 XI1.XI0.CK_EN<8> XI1.XI0.XI14<8>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<8>.MM_i_51_7 XI1.XI0.CK_EN<8> XI1.XI0.XI14<8>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<8>.MM_i_57 VDD! XI1.XI0.XI14<8>.NET_002 XI1.XI0.XI14<8>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<8>.MM_i_78 VDD! XI1.WR_ADDR_EN<8> XI1.XI0.XI14<8>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<8>.MM_i_74 XI1.XI0.XI14<8>.NET_009 XI1.XI0.XI14<8>.NET_004
+ XI1.XI0.XI14<8>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<8>.MM_i_68 XI1.XI0.XI14<8>.NET_002 XI1.XI0.XI14<8>.NET_005
+ XI1.XI0.XI14<8>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<8>.MM_i_64 XI1.XI0.XI14<8>.NET_008 XI1.XI0.XI14<8>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<8>.MM_i_84 XI1.XI0.XI14<8>.NET_004 XI1.XI0.XI14<8>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<8>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<8>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<8>.MM_i_97 XI1.XI0.XI14<8>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<8>.MM_i_103 VDD! XI1.XI0.XI14<8>.NET_000 XI1.XI0.XI14<8>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<8>.MM_i_109 XI1.XI0.CK_EN<8> XI1.XI0.XI14<8>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<8>.MM_i_109_4 XI1.XI0.CK_EN<8> XI1.XI0.XI14<8>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<7>.MM_i_0 VSS! XI1.XI0.XI14<7>.NET_002 XI1.XI0.XI14<7>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<7>.MM_i_21 VSS! XI1.WR_ADDR_EN<7> XI1.XI0.XI14<7>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<7>.MM_i_17 XI1.XI0.XI14<7>.NET_003 XI1.XI0.XI14<7>.NET_005
+ XI1.XI0.XI14<7>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<7>.MM_i_11 XI1.XI0.XI14<7>.NET_002 XI1.XI0.XI14<7>.NET_004
+ XI1.XI0.XI14<7>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<7>.MM_i_7 XI1.XI0.XI14<7>.NET_001 XI1.XI0.XI14<7>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<7>.MM_i_27 XI1.XI0.XI14<7>.NET_004 XI1.XI0.XI14<7>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<7>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<7>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<7>.MM_i_40 XI1.XI0.XI14<7>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<7>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<7>.MM_i_45 VSS! XI1.XI0.XI14<7>.NET_000 XI1.XI0.XI14<7>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<7>.MM_i_51 XI1.XI0.CK_EN<7> XI1.XI0.XI14<7>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<7>.MM_i_51_7 XI1.XI0.CK_EN<7> XI1.XI0.XI14<7>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<7>.MM_i_57 VDD! XI1.XI0.XI14<7>.NET_002 XI1.XI0.XI14<7>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<7>.MM_i_78 VDD! XI1.WR_ADDR_EN<7> XI1.XI0.XI14<7>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<7>.MM_i_74 XI1.XI0.XI14<7>.NET_009 XI1.XI0.XI14<7>.NET_004
+ XI1.XI0.XI14<7>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<7>.MM_i_68 XI1.XI0.XI14<7>.NET_002 XI1.XI0.XI14<7>.NET_005
+ XI1.XI0.XI14<7>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<7>.MM_i_64 XI1.XI0.XI14<7>.NET_008 XI1.XI0.XI14<7>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<7>.MM_i_84 XI1.XI0.XI14<7>.NET_004 XI1.XI0.XI14<7>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<7>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<7>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<7>.MM_i_97 XI1.XI0.XI14<7>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<7>.MM_i_103 VDD! XI1.XI0.XI14<7>.NET_000 XI1.XI0.XI14<7>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<7>.MM_i_109 XI1.XI0.CK_EN<7> XI1.XI0.XI14<7>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<7>.MM_i_109_4 XI1.XI0.CK_EN<7> XI1.XI0.XI14<7>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<6>.MM_i_0 VSS! XI1.XI0.XI14<6>.NET_002 XI1.XI0.XI14<6>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<6>.MM_i_21 VSS! XI1.WR_ADDR_EN<6> XI1.XI0.XI14<6>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<6>.MM_i_17 XI1.XI0.XI14<6>.NET_003 XI1.XI0.XI14<6>.NET_005
+ XI1.XI0.XI14<6>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<6>.MM_i_11 XI1.XI0.XI14<6>.NET_002 XI1.XI0.XI14<6>.NET_004
+ XI1.XI0.XI14<6>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<6>.MM_i_7 XI1.XI0.XI14<6>.NET_001 XI1.XI0.XI14<6>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<6>.MM_i_27 XI1.XI0.XI14<6>.NET_004 XI1.XI0.XI14<6>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<6>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<6>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<6>.MM_i_40 XI1.XI0.XI14<6>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<6>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<6>.MM_i_45 VSS! XI1.XI0.XI14<6>.NET_000 XI1.XI0.XI14<6>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<6>.MM_i_51 XI1.XI0.CK_EN<6> XI1.XI0.XI14<6>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<6>.MM_i_51_7 XI1.XI0.CK_EN<6> XI1.XI0.XI14<6>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<6>.MM_i_57 VDD! XI1.XI0.XI14<6>.NET_002 XI1.XI0.XI14<6>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<6>.MM_i_78 VDD! XI1.WR_ADDR_EN<6> XI1.XI0.XI14<6>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<6>.MM_i_74 XI1.XI0.XI14<6>.NET_009 XI1.XI0.XI14<6>.NET_004
+ XI1.XI0.XI14<6>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<6>.MM_i_68 XI1.XI0.XI14<6>.NET_002 XI1.XI0.XI14<6>.NET_005
+ XI1.XI0.XI14<6>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<6>.MM_i_64 XI1.XI0.XI14<6>.NET_008 XI1.XI0.XI14<6>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<6>.MM_i_84 XI1.XI0.XI14<6>.NET_004 XI1.XI0.XI14<6>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<6>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<6>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<6>.MM_i_97 XI1.XI0.XI14<6>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<6>.MM_i_103 VDD! XI1.XI0.XI14<6>.NET_000 XI1.XI0.XI14<6>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<6>.MM_i_109 XI1.XI0.CK_EN<6> XI1.XI0.XI14<6>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<6>.MM_i_109_4 XI1.XI0.CK_EN<6> XI1.XI0.XI14<6>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<5>.MM_i_0 VSS! XI1.XI0.XI14<5>.NET_002 XI1.XI0.XI14<5>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<5>.MM_i_21 VSS! XI1.WR_ADDR_EN<5> XI1.XI0.XI14<5>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<5>.MM_i_17 XI1.XI0.XI14<5>.NET_003 XI1.XI0.XI14<5>.NET_005
+ XI1.XI0.XI14<5>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<5>.MM_i_11 XI1.XI0.XI14<5>.NET_002 XI1.XI0.XI14<5>.NET_004
+ XI1.XI0.XI14<5>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<5>.MM_i_7 XI1.XI0.XI14<5>.NET_001 XI1.XI0.XI14<5>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<5>.MM_i_27 XI1.XI0.XI14<5>.NET_004 XI1.XI0.XI14<5>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<5>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<5>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<5>.MM_i_40 XI1.XI0.XI14<5>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<5>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<5>.MM_i_45 VSS! XI1.XI0.XI14<5>.NET_000 XI1.XI0.XI14<5>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<5>.MM_i_51 XI1.XI0.CK_EN<5> XI1.XI0.XI14<5>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<5>.MM_i_51_7 XI1.XI0.CK_EN<5> XI1.XI0.XI14<5>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<5>.MM_i_57 VDD! XI1.XI0.XI14<5>.NET_002 XI1.XI0.XI14<5>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<5>.MM_i_78 VDD! XI1.WR_ADDR_EN<5> XI1.XI0.XI14<5>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<5>.MM_i_74 XI1.XI0.XI14<5>.NET_009 XI1.XI0.XI14<5>.NET_004
+ XI1.XI0.XI14<5>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<5>.MM_i_68 XI1.XI0.XI14<5>.NET_002 XI1.XI0.XI14<5>.NET_005
+ XI1.XI0.XI14<5>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<5>.MM_i_64 XI1.XI0.XI14<5>.NET_008 XI1.XI0.XI14<5>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<5>.MM_i_84 XI1.XI0.XI14<5>.NET_004 XI1.XI0.XI14<5>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<5>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<5>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<5>.MM_i_97 XI1.XI0.XI14<5>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<5>.MM_i_103 VDD! XI1.XI0.XI14<5>.NET_000 XI1.XI0.XI14<5>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<5>.MM_i_109 XI1.XI0.CK_EN<5> XI1.XI0.XI14<5>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<5>.MM_i_109_4 XI1.XI0.CK_EN<5> XI1.XI0.XI14<5>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<4>.MM_i_0 VSS! XI1.XI0.XI14<4>.NET_002 XI1.XI0.XI14<4>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<4>.MM_i_21 VSS! XI1.WR_ADDR_EN<4> XI1.XI0.XI14<4>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<4>.MM_i_17 XI1.XI0.XI14<4>.NET_003 XI1.XI0.XI14<4>.NET_005
+ XI1.XI0.XI14<4>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<4>.MM_i_11 XI1.XI0.XI14<4>.NET_002 XI1.XI0.XI14<4>.NET_004
+ XI1.XI0.XI14<4>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<4>.MM_i_7 XI1.XI0.XI14<4>.NET_001 XI1.XI0.XI14<4>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<4>.MM_i_27 XI1.XI0.XI14<4>.NET_004 XI1.XI0.XI14<4>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<4>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<4>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<4>.MM_i_40 XI1.XI0.XI14<4>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<4>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<4>.MM_i_45 VSS! XI1.XI0.XI14<4>.NET_000 XI1.XI0.XI14<4>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<4>.MM_i_51 XI1.XI0.CK_EN<4> XI1.XI0.XI14<4>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<4>.MM_i_51_7 XI1.XI0.CK_EN<4> XI1.XI0.XI14<4>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<4>.MM_i_57 VDD! XI1.XI0.XI14<4>.NET_002 XI1.XI0.XI14<4>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<4>.MM_i_78 VDD! XI1.WR_ADDR_EN<4> XI1.XI0.XI14<4>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<4>.MM_i_74 XI1.XI0.XI14<4>.NET_009 XI1.XI0.XI14<4>.NET_004
+ XI1.XI0.XI14<4>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<4>.MM_i_68 XI1.XI0.XI14<4>.NET_002 XI1.XI0.XI14<4>.NET_005
+ XI1.XI0.XI14<4>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<4>.MM_i_64 XI1.XI0.XI14<4>.NET_008 XI1.XI0.XI14<4>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<4>.MM_i_84 XI1.XI0.XI14<4>.NET_004 XI1.XI0.XI14<4>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<4>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<4>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<4>.MM_i_97 XI1.XI0.XI14<4>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<4>.MM_i_103 VDD! XI1.XI0.XI14<4>.NET_000 XI1.XI0.XI14<4>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<4>.MM_i_109 XI1.XI0.CK_EN<4> XI1.XI0.XI14<4>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<4>.MM_i_109_4 XI1.XI0.CK_EN<4> XI1.XI0.XI14<4>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<3>.MM_i_0 VSS! XI1.XI0.XI14<3>.NET_002 XI1.XI0.XI14<3>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<3>.MM_i_21 VSS! XI1.WR_ADDR_EN<3> XI1.XI0.XI14<3>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<3>.MM_i_17 XI1.XI0.XI14<3>.NET_003 XI1.XI0.XI14<3>.NET_005
+ XI1.XI0.XI14<3>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<3>.MM_i_11 XI1.XI0.XI14<3>.NET_002 XI1.XI0.XI14<3>.NET_004
+ XI1.XI0.XI14<3>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<3>.MM_i_7 XI1.XI0.XI14<3>.NET_001 XI1.XI0.XI14<3>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<3>.MM_i_27 XI1.XI0.XI14<3>.NET_004 XI1.XI0.XI14<3>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<3>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<3>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<3>.MM_i_40 XI1.XI0.XI14<3>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<3>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<3>.MM_i_45 VSS! XI1.XI0.XI14<3>.NET_000 XI1.XI0.XI14<3>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<3>.MM_i_51 XI1.XI0.CK_EN<3> XI1.XI0.XI14<3>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<3>.MM_i_51_7 XI1.XI0.CK_EN<3> XI1.XI0.XI14<3>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<3>.MM_i_57 VDD! XI1.XI0.XI14<3>.NET_002 XI1.XI0.XI14<3>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<3>.MM_i_78 VDD! XI1.WR_ADDR_EN<3> XI1.XI0.XI14<3>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<3>.MM_i_74 XI1.XI0.XI14<3>.NET_009 XI1.XI0.XI14<3>.NET_004
+ XI1.XI0.XI14<3>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<3>.MM_i_68 XI1.XI0.XI14<3>.NET_002 XI1.XI0.XI14<3>.NET_005
+ XI1.XI0.XI14<3>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<3>.MM_i_64 XI1.XI0.XI14<3>.NET_008 XI1.XI0.XI14<3>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<3>.MM_i_84 XI1.XI0.XI14<3>.NET_004 XI1.XI0.XI14<3>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<3>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<3>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<3>.MM_i_97 XI1.XI0.XI14<3>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<3>.MM_i_103 VDD! XI1.XI0.XI14<3>.NET_000 XI1.XI0.XI14<3>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<3>.MM_i_109 XI1.XI0.CK_EN<3> XI1.XI0.XI14<3>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<3>.MM_i_109_4 XI1.XI0.CK_EN<3> XI1.XI0.XI14<3>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<2>.MM_i_0 VSS! XI1.XI0.XI14<2>.NET_002 XI1.XI0.XI14<2>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<2>.MM_i_21 VSS! XI1.WR_ADDR_EN<2> XI1.XI0.XI14<2>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<2>.MM_i_17 XI1.XI0.XI14<2>.NET_003 XI1.XI0.XI14<2>.NET_005
+ XI1.XI0.XI14<2>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<2>.MM_i_11 XI1.XI0.XI14<2>.NET_002 XI1.XI0.XI14<2>.NET_004
+ XI1.XI0.XI14<2>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<2>.MM_i_7 XI1.XI0.XI14<2>.NET_001 XI1.XI0.XI14<2>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<2>.MM_i_27 XI1.XI0.XI14<2>.NET_004 XI1.XI0.XI14<2>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<2>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<2>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<2>.MM_i_40 XI1.XI0.XI14<2>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<2>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<2>.MM_i_45 VSS! XI1.XI0.XI14<2>.NET_000 XI1.XI0.XI14<2>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<2>.MM_i_51 XI1.XI0.CK_EN<2> XI1.XI0.XI14<2>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<2>.MM_i_51_7 XI1.XI0.CK_EN<2> XI1.XI0.XI14<2>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<2>.MM_i_57 VDD! XI1.XI0.XI14<2>.NET_002 XI1.XI0.XI14<2>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<2>.MM_i_78 VDD! XI1.WR_ADDR_EN<2> XI1.XI0.XI14<2>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<2>.MM_i_74 XI1.XI0.XI14<2>.NET_009 XI1.XI0.XI14<2>.NET_004
+ XI1.XI0.XI14<2>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<2>.MM_i_68 XI1.XI0.XI14<2>.NET_002 XI1.XI0.XI14<2>.NET_005
+ XI1.XI0.XI14<2>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<2>.MM_i_64 XI1.XI0.XI14<2>.NET_008 XI1.XI0.XI14<2>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<2>.MM_i_84 XI1.XI0.XI14<2>.NET_004 XI1.XI0.XI14<2>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<2>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<2>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<2>.MM_i_97 XI1.XI0.XI14<2>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<2>.MM_i_103 VDD! XI1.XI0.XI14<2>.NET_000 XI1.XI0.XI14<2>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<2>.MM_i_109 XI1.XI0.CK_EN<2> XI1.XI0.XI14<2>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<2>.MM_i_109_4 XI1.XI0.CK_EN<2> XI1.XI0.XI14<2>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<1>.MM_i_0 VSS! XI1.XI0.XI14<1>.NET_002 XI1.XI0.XI14<1>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<1>.MM_i_21 VSS! XI1.WR_ADDR_EN<1> XI1.XI0.XI14<1>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<1>.MM_i_17 XI1.XI0.XI14<1>.NET_003 XI1.XI0.XI14<1>.NET_005
+ XI1.XI0.XI14<1>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<1>.MM_i_11 XI1.XI0.XI14<1>.NET_002 XI1.XI0.XI14<1>.NET_004
+ XI1.XI0.XI14<1>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<1>.MM_i_7 XI1.XI0.XI14<1>.NET_001 XI1.XI0.XI14<1>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<1>.MM_i_27 XI1.XI0.XI14<1>.NET_004 XI1.XI0.XI14<1>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<1>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<1>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<1>.MM_i_40 XI1.XI0.XI14<1>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<1>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<1>.MM_i_45 VSS! XI1.XI0.XI14<1>.NET_000 XI1.XI0.XI14<1>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<1>.MM_i_51 XI1.XI0.CK_EN<1> XI1.XI0.XI14<1>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<1>.MM_i_51_7 XI1.XI0.CK_EN<1> XI1.XI0.XI14<1>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<1>.MM_i_57 VDD! XI1.XI0.XI14<1>.NET_002 XI1.XI0.XI14<1>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<1>.MM_i_78 VDD! XI1.WR_ADDR_EN<1> XI1.XI0.XI14<1>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<1>.MM_i_74 XI1.XI0.XI14<1>.NET_009 XI1.XI0.XI14<1>.NET_004
+ XI1.XI0.XI14<1>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<1>.MM_i_68 XI1.XI0.XI14<1>.NET_002 XI1.XI0.XI14<1>.NET_005
+ XI1.XI0.XI14<1>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<1>.MM_i_64 XI1.XI0.XI14<1>.NET_008 XI1.XI0.XI14<1>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<1>.MM_i_84 XI1.XI0.XI14<1>.NET_004 XI1.XI0.XI14<1>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<1>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<1>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<1>.MM_i_97 XI1.XI0.XI14<1>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<1>.MM_i_103 VDD! XI1.XI0.XI14<1>.NET_000 XI1.XI0.XI14<1>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<1>.MM_i_109 XI1.XI0.CK_EN<1> XI1.XI0.XI14<1>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<1>.MM_i_109_4 XI1.XI0.CK_EN<1> XI1.XI0.XI14<1>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI14<0>.MM_i_0 VSS! XI1.XI0.XI14<0>.NET_002 XI1.XI0.XI14<0>.NET_000
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI14<0>.MM_i_21 VSS! XI1.WR_ADDR_EN<0> XI1.XI0.XI14<0>.NET_003 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<0>.MM_i_17 XI1.XI0.XI14<0>.NET_003 XI1.XI0.XI14<0>.NET_005
+ XI1.XI0.XI14<0>.NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.22e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI14<0>.MM_i_11 XI1.XI0.XI14<0>.NET_002 XI1.XI0.XI14<0>.NET_004
+ XI1.XI0.XI14<0>.NET_001 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=2.22e-14 AS=1.26e-14
+ PD=7e-07 PS=4.6e-07
mXI1.XI0.XI14<0>.MM_i_7 XI1.XI0.XI14<0>.NET_001 XI1.XI0.XI14<0>.NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.22e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI14<0>.MM_i_27 XI1.XI0.XI14<0>.NET_004 XI1.XI0.XI14<0>.NET_005 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.22e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI14<0>.MM_i_33 VSS! XI1.XI0.CK XI1.XI0.XI14<0>.NET_005 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.205e-14 PD=6.3e-07 PS=6.3e-07
mXI1.XI0.XI14<0>.MM_i_40 XI1.XI0.XI14<0>.NET_007 XI1.XI0.CK
+ XI1.XI0.XI14<0>.NET_006 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI14<0>.MM_i_45 VSS! XI1.XI0.XI14<0>.NET_000 XI1.XI0.XI14<0>.NET_007
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.7575e-14 AS=5.81e-14 PD=1.16e-06
+ PS=1.11e-06
mXI1.XI0.XI14<0>.MM_i_51 XI1.XI0.CK_EN<0> XI1.XI0.XI14<0>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.7575e-14 PD=6.7e-07 PS=1.16e-06
mXI1.XI0.XI14<0>.MM_i_51_7 XI1.XI0.CK_EN<0> XI1.XI0.XI14<0>.NET_006 VSS! VSS!
+ NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI14<0>.MM_i_57 VDD! XI1.XI0.XI14<0>.NET_002 XI1.XI0.XI14<0>.NET_000
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07
+ PS=8.4e-07
mXI1.XI0.XI14<0>.MM_i_78 VDD! XI1.WR_ADDR_EN<0> XI1.XI0.XI14<0>.NET_009 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<0>.MM_i_74 XI1.XI0.XI14<0>.NET_009 XI1.XI0.XI14<0>.NET_004
+ XI1.XI0.XI14<0>.NET_002 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.06e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI14<0>.MM_i_68 XI1.XI0.XI14<0>.NET_002 XI1.XI0.XI14<0>.NET_005
+ XI1.XI0.XI14<0>.NET_008 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=3.06e-14 AS=1.26e-14
+ PD=9.1e-07 PS=4.6e-07
mXI1.XI0.XI14<0>.MM_i_64 XI1.XI0.XI14<0>.NET_008 XI1.XI0.XI14<0>.NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.1725e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI14<0>.MM_i_84 XI1.XI0.XI14<0>.NET_004 XI1.XI0.XI14<0>.NET_005 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=3.1725e-14 PD=9.9e-07
+ PS=9.1e-07
mXI1.XI0.XI14<0>.MM_i_90 VDD! XI1.XI0.CK XI1.XI0.XI14<0>.NET_005 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.06e-06
mXI1.XI0.XI14<0>.MM_i_97 XI1.XI0.XI14<0>.NET_006 XI1.XI0.CK VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI14<0>.MM_i_103 VDD! XI1.XI0.XI14<0>.NET_000 XI1.XI0.XI14<0>.NET_006
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=1.0395e-13 AS=8.82e-14 PD=1.59e-06
+ PS=1.54e-06
mXI1.XI0.XI14<0>.MM_i_109 XI1.XI0.CK_EN<0> XI1.XI0.XI14<0>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.0395e-13 PD=1.54e-06 PS=1.59e-06
mXI1.XI0.XI14<0>.MM_i_109_4 XI1.XI0.CK_EN<0> XI1.XI0.XI14<0>.NET_006 VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI1<12>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_41_11 REG_DATA_12<3> XI1.XI0.XI1<12>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<3>.MM_i_7 XI1.XI0.XI1<12>.XI7<3>.NET_001
+ XI1.XI0.XI1<12>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_13 XI1.XI0.XI1<12>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_18 XI1.XI0.XI1<12>.XI7<3>.NET_003
+ XI1.XI0.XI1<12>.XI7<3>.NET_001 XI1.XI0.XI1<12>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_24 XI1.XI0.XI1<12>.XI7<3>.NET_004
+ XI1.XI0.XI1<12>.XI7<3>.NET_000 XI1.XI0.XI1<12>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<3>.NET_005
+ XI1.XI0.XI1<12>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<3>.NET_003
+ XI1.XI0.XI1<12>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_89_4 REG_DATA_12<3> XI1.XI0.XI1<12>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<3>.MM_i_55 XI1.XI0.XI1<12>.XI7<3>.NET_001
+ XI1.XI0.XI1<12>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_61 XI1.XI0.XI1<12>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_66 XI1.XI0.XI1<12>.XI7<3>.NET_003
+ XI1.XI0.XI1<12>.XI7<3>.NET_000 XI1.XI0.XI1<12>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_72 XI1.XI0.XI1<12>.XI7<3>.NET_007
+ XI1.XI0.XI1<12>.XI7<3>.NET_001 XI1.XI0.XI1<12>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<3>.NET_005
+ XI1.XI0.XI1<12>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<3>.NET_003
+ XI1.XI0.XI1<12>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_41_11 REG_DATA_12<2> XI1.XI0.XI1<12>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<2>.MM_i_7 XI1.XI0.XI1<12>.XI7<2>.NET_001
+ XI1.XI0.XI1<12>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_13 XI1.XI0.XI1<12>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_18 XI1.XI0.XI1<12>.XI7<2>.NET_003
+ XI1.XI0.XI1<12>.XI7<2>.NET_001 XI1.XI0.XI1<12>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_24 XI1.XI0.XI1<12>.XI7<2>.NET_004
+ XI1.XI0.XI1<12>.XI7<2>.NET_000 XI1.XI0.XI1<12>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<2>.NET_005
+ XI1.XI0.XI1<12>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<2>.NET_003
+ XI1.XI0.XI1<12>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_89_4 REG_DATA_12<2> XI1.XI0.XI1<12>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<2>.MM_i_55 XI1.XI0.XI1<12>.XI7<2>.NET_001
+ XI1.XI0.XI1<12>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_61 XI1.XI0.XI1<12>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_66 XI1.XI0.XI1<12>.XI7<2>.NET_003
+ XI1.XI0.XI1<12>.XI7<2>.NET_000 XI1.XI0.XI1<12>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_72 XI1.XI0.XI1<12>.XI7<2>.NET_007
+ XI1.XI0.XI1<12>.XI7<2>.NET_001 XI1.XI0.XI1<12>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<2>.NET_005
+ XI1.XI0.XI1<12>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<2>.NET_003
+ XI1.XI0.XI1<12>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_41_11 REG_DATA_12<1> XI1.XI0.XI1<12>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<1>.MM_i_7 XI1.XI0.XI1<12>.XI7<1>.NET_001
+ XI1.XI0.XI1<12>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_13 XI1.XI0.XI1<12>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_18 XI1.XI0.XI1<12>.XI7<1>.NET_003
+ XI1.XI0.XI1<12>.XI7<1>.NET_001 XI1.XI0.XI1<12>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_24 XI1.XI0.XI1<12>.XI7<1>.NET_004
+ XI1.XI0.XI1<12>.XI7<1>.NET_000 XI1.XI0.XI1<12>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<1>.NET_005
+ XI1.XI0.XI1<12>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<1>.NET_003
+ XI1.XI0.XI1<12>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_89_4 REG_DATA_12<1> XI1.XI0.XI1<12>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<1>.MM_i_55 XI1.XI0.XI1<12>.XI7<1>.NET_001
+ XI1.XI0.XI1<12>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_61 XI1.XI0.XI1<12>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_66 XI1.XI0.XI1<12>.XI7<1>.NET_003
+ XI1.XI0.XI1<12>.XI7<1>.NET_000 XI1.XI0.XI1<12>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_72 XI1.XI0.XI1<12>.XI7<1>.NET_007
+ XI1.XI0.XI1<12>.XI7<1>.NET_001 XI1.XI0.XI1<12>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<1>.NET_005
+ XI1.XI0.XI1<12>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<1>.NET_003
+ XI1.XI0.XI1<12>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_41_11 REG_DATA_12<0> XI1.XI0.XI1<12>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<0>.MM_i_7 XI1.XI0.XI1<12>.XI7<0>.NET_001
+ XI1.XI0.XI1<12>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_13 XI1.XI0.XI1<12>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_18 XI1.XI0.XI1<12>.XI7<0>.NET_003
+ XI1.XI0.XI1<12>.XI7<0>.NET_001 XI1.XI0.XI1<12>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_24 XI1.XI0.XI1<12>.XI7<0>.NET_004
+ XI1.XI0.XI1<12>.XI7<0>.NET_000 XI1.XI0.XI1<12>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<0>.NET_005
+ XI1.XI0.XI1<12>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<0>.NET_003
+ XI1.XI0.XI1<12>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_89_4 REG_DATA_12<0> XI1.XI0.XI1<12>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<0>.MM_i_55 XI1.XI0.XI1<12>.XI7<0>.NET_001
+ XI1.XI0.XI1<12>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_61 XI1.XI0.XI1<12>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_66 XI1.XI0.XI1<12>.XI7<0>.NET_003
+ XI1.XI0.XI1<12>.XI7<0>.NET_000 XI1.XI0.XI1<12>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_72 XI1.XI0.XI1<12>.XI7<0>.NET_007
+ XI1.XI0.XI1<12>.XI7<0>.NET_001 XI1.XI0.XI1<12>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<0>.NET_005
+ XI1.XI0.XI1<12>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<0>.NET_003
+ XI1.XI0.XI1<12>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_41_11 REG_DATA_12<7> XI1.XI0.XI1<12>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<7>.MM_i_7 XI1.XI0.XI1<12>.XI7<7>.NET_001
+ XI1.XI0.XI1<12>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_13 XI1.XI0.XI1<12>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_18 XI1.XI0.XI1<12>.XI7<7>.NET_003
+ XI1.XI0.XI1<12>.XI7<7>.NET_001 XI1.XI0.XI1<12>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_24 XI1.XI0.XI1<12>.XI7<7>.NET_004
+ XI1.XI0.XI1<12>.XI7<7>.NET_000 XI1.XI0.XI1<12>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<7>.NET_005
+ XI1.XI0.XI1<12>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<7>.NET_003
+ XI1.XI0.XI1<12>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_89_4 REG_DATA_12<7> XI1.XI0.XI1<12>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<7>.MM_i_55 XI1.XI0.XI1<12>.XI7<7>.NET_001
+ XI1.XI0.XI1<12>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_61 XI1.XI0.XI1<12>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_66 XI1.XI0.XI1<12>.XI7<7>.NET_003
+ XI1.XI0.XI1<12>.XI7<7>.NET_000 XI1.XI0.XI1<12>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_72 XI1.XI0.XI1<12>.XI7<7>.NET_007
+ XI1.XI0.XI1<12>.XI7<7>.NET_001 XI1.XI0.XI1<12>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<7>.NET_005
+ XI1.XI0.XI1<12>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<7>.NET_003
+ XI1.XI0.XI1<12>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_41_11 REG_DATA_12<6> XI1.XI0.XI1<12>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<6>.MM_i_7 XI1.XI0.XI1<12>.XI7<6>.NET_001
+ XI1.XI0.XI1<12>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_13 XI1.XI0.XI1<12>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_18 XI1.XI0.XI1<12>.XI7<6>.NET_003
+ XI1.XI0.XI1<12>.XI7<6>.NET_001 XI1.XI0.XI1<12>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_24 XI1.XI0.XI1<12>.XI7<6>.NET_004
+ XI1.XI0.XI1<12>.XI7<6>.NET_000 XI1.XI0.XI1<12>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<6>.NET_005
+ XI1.XI0.XI1<12>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<6>.NET_003
+ XI1.XI0.XI1<12>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_89_4 REG_DATA_12<6> XI1.XI0.XI1<12>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<6>.MM_i_55 XI1.XI0.XI1<12>.XI7<6>.NET_001
+ XI1.XI0.XI1<12>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_61 XI1.XI0.XI1<12>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_66 XI1.XI0.XI1<12>.XI7<6>.NET_003
+ XI1.XI0.XI1<12>.XI7<6>.NET_000 XI1.XI0.XI1<12>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_72 XI1.XI0.XI1<12>.XI7<6>.NET_007
+ XI1.XI0.XI1<12>.XI7<6>.NET_001 XI1.XI0.XI1<12>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<6>.NET_005
+ XI1.XI0.XI1<12>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<6>.NET_003
+ XI1.XI0.XI1<12>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_41_11 REG_DATA_12<5> XI1.XI0.XI1<12>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<5>.MM_i_7 XI1.XI0.XI1<12>.XI7<5>.NET_001
+ XI1.XI0.XI1<12>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_13 XI1.XI0.XI1<12>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_18 XI1.XI0.XI1<12>.XI7<5>.NET_003
+ XI1.XI0.XI1<12>.XI7<5>.NET_001 XI1.XI0.XI1<12>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_24 XI1.XI0.XI1<12>.XI7<5>.NET_004
+ XI1.XI0.XI1<12>.XI7<5>.NET_000 XI1.XI0.XI1<12>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<5>.NET_005
+ XI1.XI0.XI1<12>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<5>.NET_003
+ XI1.XI0.XI1<12>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_89_4 REG_DATA_12<5> XI1.XI0.XI1<12>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<5>.MM_i_55 XI1.XI0.XI1<12>.XI7<5>.NET_001
+ XI1.XI0.XI1<12>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_61 XI1.XI0.XI1<12>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_66 XI1.XI0.XI1<12>.XI7<5>.NET_003
+ XI1.XI0.XI1<12>.XI7<5>.NET_000 XI1.XI0.XI1<12>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_72 XI1.XI0.XI1<12>.XI7<5>.NET_007
+ XI1.XI0.XI1<12>.XI7<5>.NET_001 XI1.XI0.XI1<12>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<5>.NET_005
+ XI1.XI0.XI1<12>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<5>.NET_003
+ XI1.XI0.XI1<12>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_41_11 REG_DATA_12<4> XI1.XI0.XI1<12>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<4>.MM_i_7 XI1.XI0.XI1<12>.XI7<4>.NET_001
+ XI1.XI0.XI1<12>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_13 XI1.XI0.XI1<12>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_18 XI1.XI0.XI1<12>.XI7<4>.NET_003
+ XI1.XI0.XI1<12>.XI7<4>.NET_001 XI1.XI0.XI1<12>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_24 XI1.XI0.XI1<12>.XI7<4>.NET_004
+ XI1.XI0.XI1<12>.XI7<4>.NET_000 XI1.XI0.XI1<12>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<4>.NET_005
+ XI1.XI0.XI1<12>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<4>.NET_003
+ XI1.XI0.XI1<12>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_89_4 REG_DATA_12<4> XI1.XI0.XI1<12>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<4>.MM_i_55 XI1.XI0.XI1<12>.XI7<4>.NET_001
+ XI1.XI0.XI1<12>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_61 XI1.XI0.XI1<12>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_66 XI1.XI0.XI1<12>.XI7<4>.NET_003
+ XI1.XI0.XI1<12>.XI7<4>.NET_000 XI1.XI0.XI1<12>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_72 XI1.XI0.XI1<12>.XI7<4>.NET_007
+ XI1.XI0.XI1<12>.XI7<4>.NET_001 XI1.XI0.XI1<12>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<4>.NET_005
+ XI1.XI0.XI1<12>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<4>.NET_003
+ XI1.XI0.XI1<12>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_41_11 REG_DATA_12<11>
+ XI1.XI0.XI1<12>.XI7<11>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<11>.MM_i_7 XI1.XI0.XI1<12>.XI7<11>.NET_001
+ XI1.XI0.XI1<12>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_13 XI1.XI0.XI1<12>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_18 XI1.XI0.XI1<12>.XI7<11>.NET_003
+ XI1.XI0.XI1<12>.XI7<11>.NET_001 XI1.XI0.XI1<12>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_24 XI1.XI0.XI1<12>.XI7<11>.NET_004
+ XI1.XI0.XI1<12>.XI7<11>.NET_000 XI1.XI0.XI1<12>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<11>.NET_005
+ XI1.XI0.XI1<12>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<11>.NET_003
+ XI1.XI0.XI1<12>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_89_4 REG_DATA_12<11>
+ XI1.XI0.XI1<12>.XI7<11>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<11>.MM_i_55 XI1.XI0.XI1<12>.XI7<11>.NET_001
+ XI1.XI0.XI1<12>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_61 XI1.XI0.XI1<12>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_66 XI1.XI0.XI1<12>.XI7<11>.NET_003
+ XI1.XI0.XI1<12>.XI7<11>.NET_000 XI1.XI0.XI1<12>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_72 XI1.XI0.XI1<12>.XI7<11>.NET_007
+ XI1.XI0.XI1<12>.XI7<11>.NET_001 XI1.XI0.XI1<12>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<11>.NET_005
+ XI1.XI0.XI1<12>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<11>.NET_003
+ XI1.XI0.XI1<12>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_41_11 REG_DATA_12<10>
+ XI1.XI0.XI1<12>.XI7<10>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<10>.MM_i_7 XI1.XI0.XI1<12>.XI7<10>.NET_001
+ XI1.XI0.XI1<12>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_13 XI1.XI0.XI1<12>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_18 XI1.XI0.XI1<12>.XI7<10>.NET_003
+ XI1.XI0.XI1<12>.XI7<10>.NET_001 XI1.XI0.XI1<12>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_24 XI1.XI0.XI1<12>.XI7<10>.NET_004
+ XI1.XI0.XI1<12>.XI7<10>.NET_000 XI1.XI0.XI1<12>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<10>.NET_005
+ XI1.XI0.XI1<12>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<10>.NET_003
+ XI1.XI0.XI1<12>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_89_4 REG_DATA_12<10>
+ XI1.XI0.XI1<12>.XI7<10>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<10>.MM_i_55 XI1.XI0.XI1<12>.XI7<10>.NET_001
+ XI1.XI0.XI1<12>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_61 XI1.XI0.XI1<12>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_66 XI1.XI0.XI1<12>.XI7<10>.NET_003
+ XI1.XI0.XI1<12>.XI7<10>.NET_000 XI1.XI0.XI1<12>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_72 XI1.XI0.XI1<12>.XI7<10>.NET_007
+ XI1.XI0.XI1<12>.XI7<10>.NET_001 XI1.XI0.XI1<12>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<10>.NET_005
+ XI1.XI0.XI1<12>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<10>.NET_003
+ XI1.XI0.XI1<12>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_41_11 REG_DATA_12<9> XI1.XI0.XI1<12>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<9>.MM_i_7 XI1.XI0.XI1<12>.XI7<9>.NET_001
+ XI1.XI0.XI1<12>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_13 XI1.XI0.XI1<12>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_18 XI1.XI0.XI1<12>.XI7<9>.NET_003
+ XI1.XI0.XI1<12>.XI7<9>.NET_001 XI1.XI0.XI1<12>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_24 XI1.XI0.XI1<12>.XI7<9>.NET_004
+ XI1.XI0.XI1<12>.XI7<9>.NET_000 XI1.XI0.XI1<12>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<9>.NET_005
+ XI1.XI0.XI1<12>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<9>.NET_003
+ XI1.XI0.XI1<12>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_89_4 REG_DATA_12<9> XI1.XI0.XI1<12>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<9>.MM_i_55 XI1.XI0.XI1<12>.XI7<9>.NET_001
+ XI1.XI0.XI1<12>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_61 XI1.XI0.XI1<12>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_66 XI1.XI0.XI1<12>.XI7<9>.NET_003
+ XI1.XI0.XI1<12>.XI7<9>.NET_000 XI1.XI0.XI1<12>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_72 XI1.XI0.XI1<12>.XI7<9>.NET_007
+ XI1.XI0.XI1<12>.XI7<9>.NET_001 XI1.XI0.XI1<12>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<9>.NET_005
+ XI1.XI0.XI1<12>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<9>.NET_003
+ XI1.XI0.XI1<12>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_41_11 REG_DATA_12<8> XI1.XI0.XI1<12>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<8>.MM_i_7 XI1.XI0.XI1<12>.XI7<8>.NET_001
+ XI1.XI0.XI1<12>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_13 XI1.XI0.XI1<12>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_18 XI1.XI0.XI1<12>.XI7<8>.NET_003
+ XI1.XI0.XI1<12>.XI7<8>.NET_001 XI1.XI0.XI1<12>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_24 XI1.XI0.XI1<12>.XI7<8>.NET_004
+ XI1.XI0.XI1<12>.XI7<8>.NET_000 XI1.XI0.XI1<12>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<8>.NET_005
+ XI1.XI0.XI1<12>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<8>.NET_003
+ XI1.XI0.XI1<12>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_89_4 REG_DATA_12<8> XI1.XI0.XI1<12>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<8>.MM_i_55 XI1.XI0.XI1<12>.XI7<8>.NET_001
+ XI1.XI0.XI1<12>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_61 XI1.XI0.XI1<12>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_66 XI1.XI0.XI1<12>.XI7<8>.NET_003
+ XI1.XI0.XI1<12>.XI7<8>.NET_000 XI1.XI0.XI1<12>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_72 XI1.XI0.XI1<12>.XI7<8>.NET_007
+ XI1.XI0.XI1<12>.XI7<8>.NET_001 XI1.XI0.XI1<12>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<8>.NET_005
+ XI1.XI0.XI1<12>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<8>.NET_003
+ XI1.XI0.XI1<12>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_41_11 REG_DATA_12<15>
+ XI1.XI0.XI1<12>.XI7<15>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<15>.MM_i_7 XI1.XI0.XI1<12>.XI7<15>.NET_001
+ XI1.XI0.XI1<12>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_13 XI1.XI0.XI1<12>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_18 XI1.XI0.XI1<12>.XI7<15>.NET_003
+ XI1.XI0.XI1<12>.XI7<15>.NET_001 XI1.XI0.XI1<12>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_24 XI1.XI0.XI1<12>.XI7<15>.NET_004
+ XI1.XI0.XI1<12>.XI7<15>.NET_000 XI1.XI0.XI1<12>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<15>.NET_005
+ XI1.XI0.XI1<12>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<15>.NET_003
+ XI1.XI0.XI1<12>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_89_4 REG_DATA_12<15>
+ XI1.XI0.XI1<12>.XI7<15>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<15>.MM_i_55 XI1.XI0.XI1<12>.XI7<15>.NET_001
+ XI1.XI0.XI1<12>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_61 XI1.XI0.XI1<12>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_66 XI1.XI0.XI1<12>.XI7<15>.NET_003
+ XI1.XI0.XI1<12>.XI7<15>.NET_000 XI1.XI0.XI1<12>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_72 XI1.XI0.XI1<12>.XI7<15>.NET_007
+ XI1.XI0.XI1<12>.XI7<15>.NET_001 XI1.XI0.XI1<12>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<15>.NET_005
+ XI1.XI0.XI1<12>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<15>.NET_003
+ XI1.XI0.XI1<12>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_41_11 REG_DATA_12<14>
+ XI1.XI0.XI1<12>.XI7<14>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<14>.MM_i_7 XI1.XI0.XI1<12>.XI7<14>.NET_001
+ XI1.XI0.XI1<12>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_13 XI1.XI0.XI1<12>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_18 XI1.XI0.XI1<12>.XI7<14>.NET_003
+ XI1.XI0.XI1<12>.XI7<14>.NET_001 XI1.XI0.XI1<12>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_24 XI1.XI0.XI1<12>.XI7<14>.NET_004
+ XI1.XI0.XI1<12>.XI7<14>.NET_000 XI1.XI0.XI1<12>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<14>.NET_005
+ XI1.XI0.XI1<12>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<14>.NET_003
+ XI1.XI0.XI1<12>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_89_4 REG_DATA_12<14>
+ XI1.XI0.XI1<12>.XI7<14>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<14>.MM_i_55 XI1.XI0.XI1<12>.XI7<14>.NET_001
+ XI1.XI0.XI1<12>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_61 XI1.XI0.XI1<12>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_66 XI1.XI0.XI1<12>.XI7<14>.NET_003
+ XI1.XI0.XI1<12>.XI7<14>.NET_000 XI1.XI0.XI1<12>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_72 XI1.XI0.XI1<12>.XI7<14>.NET_007
+ XI1.XI0.XI1<12>.XI7<14>.NET_001 XI1.XI0.XI1<12>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<14>.NET_005
+ XI1.XI0.XI1<12>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<14>.NET_003
+ XI1.XI0.XI1<12>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_41_11 REG_DATA_12<13>
+ XI1.XI0.XI1<12>.XI7<13>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<13>.MM_i_7 XI1.XI0.XI1<12>.XI7<13>.NET_001
+ XI1.XI0.XI1<12>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_13 XI1.XI0.XI1<12>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_18 XI1.XI0.XI1<12>.XI7<13>.NET_003
+ XI1.XI0.XI1<12>.XI7<13>.NET_001 XI1.XI0.XI1<12>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_24 XI1.XI0.XI1<12>.XI7<13>.NET_004
+ XI1.XI0.XI1<12>.XI7<13>.NET_000 XI1.XI0.XI1<12>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<13>.NET_005
+ XI1.XI0.XI1<12>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<13>.NET_003
+ XI1.XI0.XI1<12>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_89_4 REG_DATA_12<13>
+ XI1.XI0.XI1<12>.XI7<13>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<13>.MM_i_55 XI1.XI0.XI1<12>.XI7<13>.NET_001
+ XI1.XI0.XI1<12>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_61 XI1.XI0.XI1<12>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_66 XI1.XI0.XI1<12>.XI7<13>.NET_003
+ XI1.XI0.XI1<12>.XI7<13>.NET_000 XI1.XI0.XI1<12>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_72 XI1.XI0.XI1<12>.XI7<13>.NET_007
+ XI1.XI0.XI1<12>.XI7<13>.NET_001 XI1.XI0.XI1<12>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<13>.NET_005
+ XI1.XI0.XI1<12>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<13>.NET_003
+ XI1.XI0.XI1<12>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_41_11 REG_DATA_12<12>
+ XI1.XI0.XI1<12>.XI7<12>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<12>.XI7<12>.MM_i_7 XI1.XI0.XI1<12>.XI7<12>.NET_001
+ XI1.XI0.XI1<12>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_13 XI1.XI0.XI1<12>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_18 XI1.XI0.XI1<12>.XI7<12>.NET_003
+ XI1.XI0.XI1<12>.XI7<12>.NET_001 XI1.XI0.XI1<12>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_24 XI1.XI0.XI1<12>.XI7<12>.NET_004
+ XI1.XI0.XI1<12>.XI7<12>.NET_000 XI1.XI0.XI1<12>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<12>.XI7<12>.NET_005
+ XI1.XI0.XI1<12>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<12>.XI7<12>.NET_003
+ XI1.XI0.XI1<12>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<12>
+ XI1.XI0.XI1<12>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_89_4 REG_DATA_12<12>
+ XI1.XI0.XI1<12>.XI7<12>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<12>.XI7<12>.MM_i_55 XI1.XI0.XI1<12>.XI7<12>.NET_001
+ XI1.XI0.XI1<12>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_61 XI1.XI0.XI1<12>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_66 XI1.XI0.XI1<12>.XI7<12>.NET_003
+ XI1.XI0.XI1<12>.XI7<12>.NET_000 XI1.XI0.XI1<12>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_72 XI1.XI0.XI1<12>.XI7<12>.NET_007
+ XI1.XI0.XI1<12>.XI7<12>.NET_001 XI1.XI0.XI1<12>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<12>.XI7<12>.NET_005
+ XI1.XI0.XI1<12>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<12>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<12>.XI7<12>.NET_003
+ XI1.XI0.XI1<12>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_41_11 REG_DATA_11<3> XI1.XI0.XI1<11>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<3>.MM_i_7 XI1.XI0.XI1<11>.XI7<3>.NET_001
+ XI1.XI0.XI1<11>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_13 XI1.XI0.XI1<11>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_18 XI1.XI0.XI1<11>.XI7<3>.NET_003
+ XI1.XI0.XI1<11>.XI7<3>.NET_001 XI1.XI0.XI1<11>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_24 XI1.XI0.XI1<11>.XI7<3>.NET_004
+ XI1.XI0.XI1<11>.XI7<3>.NET_000 XI1.XI0.XI1<11>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<3>.NET_005
+ XI1.XI0.XI1<11>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<3>.NET_003
+ XI1.XI0.XI1<11>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_89_4 REG_DATA_11<3> XI1.XI0.XI1<11>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<3>.MM_i_55 XI1.XI0.XI1<11>.XI7<3>.NET_001
+ XI1.XI0.XI1<11>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_61 XI1.XI0.XI1<11>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_66 XI1.XI0.XI1<11>.XI7<3>.NET_003
+ XI1.XI0.XI1<11>.XI7<3>.NET_000 XI1.XI0.XI1<11>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_72 XI1.XI0.XI1<11>.XI7<3>.NET_007
+ XI1.XI0.XI1<11>.XI7<3>.NET_001 XI1.XI0.XI1<11>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<3>.NET_005
+ XI1.XI0.XI1<11>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<3>.NET_003
+ XI1.XI0.XI1<11>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_41_11 REG_DATA_11<2> XI1.XI0.XI1<11>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<2>.MM_i_7 XI1.XI0.XI1<11>.XI7<2>.NET_001
+ XI1.XI0.XI1<11>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_13 XI1.XI0.XI1<11>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_18 XI1.XI0.XI1<11>.XI7<2>.NET_003
+ XI1.XI0.XI1<11>.XI7<2>.NET_001 XI1.XI0.XI1<11>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_24 XI1.XI0.XI1<11>.XI7<2>.NET_004
+ XI1.XI0.XI1<11>.XI7<2>.NET_000 XI1.XI0.XI1<11>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<2>.NET_005
+ XI1.XI0.XI1<11>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<2>.NET_003
+ XI1.XI0.XI1<11>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_89_4 REG_DATA_11<2> XI1.XI0.XI1<11>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<2>.MM_i_55 XI1.XI0.XI1<11>.XI7<2>.NET_001
+ XI1.XI0.XI1<11>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_61 XI1.XI0.XI1<11>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_66 XI1.XI0.XI1<11>.XI7<2>.NET_003
+ XI1.XI0.XI1<11>.XI7<2>.NET_000 XI1.XI0.XI1<11>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_72 XI1.XI0.XI1<11>.XI7<2>.NET_007
+ XI1.XI0.XI1<11>.XI7<2>.NET_001 XI1.XI0.XI1<11>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<2>.NET_005
+ XI1.XI0.XI1<11>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<2>.NET_003
+ XI1.XI0.XI1<11>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_41_11 REG_DATA_11<1> XI1.XI0.XI1<11>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<1>.MM_i_7 XI1.XI0.XI1<11>.XI7<1>.NET_001
+ XI1.XI0.XI1<11>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_13 XI1.XI0.XI1<11>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_18 XI1.XI0.XI1<11>.XI7<1>.NET_003
+ XI1.XI0.XI1<11>.XI7<1>.NET_001 XI1.XI0.XI1<11>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_24 XI1.XI0.XI1<11>.XI7<1>.NET_004
+ XI1.XI0.XI1<11>.XI7<1>.NET_000 XI1.XI0.XI1<11>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<1>.NET_005
+ XI1.XI0.XI1<11>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<1>.NET_003
+ XI1.XI0.XI1<11>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_89_4 REG_DATA_11<1> XI1.XI0.XI1<11>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<1>.MM_i_55 XI1.XI0.XI1<11>.XI7<1>.NET_001
+ XI1.XI0.XI1<11>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_61 XI1.XI0.XI1<11>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_66 XI1.XI0.XI1<11>.XI7<1>.NET_003
+ XI1.XI0.XI1<11>.XI7<1>.NET_000 XI1.XI0.XI1<11>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_72 XI1.XI0.XI1<11>.XI7<1>.NET_007
+ XI1.XI0.XI1<11>.XI7<1>.NET_001 XI1.XI0.XI1<11>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<1>.NET_005
+ XI1.XI0.XI1<11>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<1>.NET_003
+ XI1.XI0.XI1<11>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_41_11 REG_DATA_11<0> XI1.XI0.XI1<11>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<0>.MM_i_7 XI1.XI0.XI1<11>.XI7<0>.NET_001
+ XI1.XI0.XI1<11>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_13 XI1.XI0.XI1<11>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_18 XI1.XI0.XI1<11>.XI7<0>.NET_003
+ XI1.XI0.XI1<11>.XI7<0>.NET_001 XI1.XI0.XI1<11>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_24 XI1.XI0.XI1<11>.XI7<0>.NET_004
+ XI1.XI0.XI1<11>.XI7<0>.NET_000 XI1.XI0.XI1<11>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<0>.NET_005
+ XI1.XI0.XI1<11>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<0>.NET_003
+ XI1.XI0.XI1<11>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_89_4 REG_DATA_11<0> XI1.XI0.XI1<11>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<0>.MM_i_55 XI1.XI0.XI1<11>.XI7<0>.NET_001
+ XI1.XI0.XI1<11>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_61 XI1.XI0.XI1<11>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_66 XI1.XI0.XI1<11>.XI7<0>.NET_003
+ XI1.XI0.XI1<11>.XI7<0>.NET_000 XI1.XI0.XI1<11>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_72 XI1.XI0.XI1<11>.XI7<0>.NET_007
+ XI1.XI0.XI1<11>.XI7<0>.NET_001 XI1.XI0.XI1<11>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<0>.NET_005
+ XI1.XI0.XI1<11>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<0>.NET_003
+ XI1.XI0.XI1<11>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_41_11 REG_DATA_11<7> XI1.XI0.XI1<11>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<7>.MM_i_7 XI1.XI0.XI1<11>.XI7<7>.NET_001
+ XI1.XI0.XI1<11>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_13 XI1.XI0.XI1<11>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_18 XI1.XI0.XI1<11>.XI7<7>.NET_003
+ XI1.XI0.XI1<11>.XI7<7>.NET_001 XI1.XI0.XI1<11>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_24 XI1.XI0.XI1<11>.XI7<7>.NET_004
+ XI1.XI0.XI1<11>.XI7<7>.NET_000 XI1.XI0.XI1<11>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<7>.NET_005
+ XI1.XI0.XI1<11>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<7>.NET_003
+ XI1.XI0.XI1<11>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_89_4 REG_DATA_11<7> XI1.XI0.XI1<11>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<7>.MM_i_55 XI1.XI0.XI1<11>.XI7<7>.NET_001
+ XI1.XI0.XI1<11>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_61 XI1.XI0.XI1<11>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_66 XI1.XI0.XI1<11>.XI7<7>.NET_003
+ XI1.XI0.XI1<11>.XI7<7>.NET_000 XI1.XI0.XI1<11>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_72 XI1.XI0.XI1<11>.XI7<7>.NET_007
+ XI1.XI0.XI1<11>.XI7<7>.NET_001 XI1.XI0.XI1<11>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<7>.NET_005
+ XI1.XI0.XI1<11>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<7>.NET_003
+ XI1.XI0.XI1<11>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_41_11 REG_DATA_11<6> XI1.XI0.XI1<11>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<6>.MM_i_7 XI1.XI0.XI1<11>.XI7<6>.NET_001
+ XI1.XI0.XI1<11>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_13 XI1.XI0.XI1<11>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_18 XI1.XI0.XI1<11>.XI7<6>.NET_003
+ XI1.XI0.XI1<11>.XI7<6>.NET_001 XI1.XI0.XI1<11>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_24 XI1.XI0.XI1<11>.XI7<6>.NET_004
+ XI1.XI0.XI1<11>.XI7<6>.NET_000 XI1.XI0.XI1<11>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<6>.NET_005
+ XI1.XI0.XI1<11>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<6>.NET_003
+ XI1.XI0.XI1<11>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_89_4 REG_DATA_11<6> XI1.XI0.XI1<11>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<6>.MM_i_55 XI1.XI0.XI1<11>.XI7<6>.NET_001
+ XI1.XI0.XI1<11>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_61 XI1.XI0.XI1<11>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_66 XI1.XI0.XI1<11>.XI7<6>.NET_003
+ XI1.XI0.XI1<11>.XI7<6>.NET_000 XI1.XI0.XI1<11>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_72 XI1.XI0.XI1<11>.XI7<6>.NET_007
+ XI1.XI0.XI1<11>.XI7<6>.NET_001 XI1.XI0.XI1<11>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<6>.NET_005
+ XI1.XI0.XI1<11>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<6>.NET_003
+ XI1.XI0.XI1<11>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_41_11 REG_DATA_11<5> XI1.XI0.XI1<11>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<5>.MM_i_7 XI1.XI0.XI1<11>.XI7<5>.NET_001
+ XI1.XI0.XI1<11>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_13 XI1.XI0.XI1<11>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_18 XI1.XI0.XI1<11>.XI7<5>.NET_003
+ XI1.XI0.XI1<11>.XI7<5>.NET_001 XI1.XI0.XI1<11>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_24 XI1.XI0.XI1<11>.XI7<5>.NET_004
+ XI1.XI0.XI1<11>.XI7<5>.NET_000 XI1.XI0.XI1<11>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<5>.NET_005
+ XI1.XI0.XI1<11>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<5>.NET_003
+ XI1.XI0.XI1<11>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_89_4 REG_DATA_11<5> XI1.XI0.XI1<11>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<5>.MM_i_55 XI1.XI0.XI1<11>.XI7<5>.NET_001
+ XI1.XI0.XI1<11>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_61 XI1.XI0.XI1<11>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_66 XI1.XI0.XI1<11>.XI7<5>.NET_003
+ XI1.XI0.XI1<11>.XI7<5>.NET_000 XI1.XI0.XI1<11>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_72 XI1.XI0.XI1<11>.XI7<5>.NET_007
+ XI1.XI0.XI1<11>.XI7<5>.NET_001 XI1.XI0.XI1<11>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<5>.NET_005
+ XI1.XI0.XI1<11>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<5>.NET_003
+ XI1.XI0.XI1<11>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_41_11 REG_DATA_11<4> XI1.XI0.XI1<11>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<4>.MM_i_7 XI1.XI0.XI1<11>.XI7<4>.NET_001
+ XI1.XI0.XI1<11>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_13 XI1.XI0.XI1<11>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_18 XI1.XI0.XI1<11>.XI7<4>.NET_003
+ XI1.XI0.XI1<11>.XI7<4>.NET_001 XI1.XI0.XI1<11>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_24 XI1.XI0.XI1<11>.XI7<4>.NET_004
+ XI1.XI0.XI1<11>.XI7<4>.NET_000 XI1.XI0.XI1<11>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<4>.NET_005
+ XI1.XI0.XI1<11>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<4>.NET_003
+ XI1.XI0.XI1<11>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_89_4 REG_DATA_11<4> XI1.XI0.XI1<11>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<4>.MM_i_55 XI1.XI0.XI1<11>.XI7<4>.NET_001
+ XI1.XI0.XI1<11>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_61 XI1.XI0.XI1<11>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_66 XI1.XI0.XI1<11>.XI7<4>.NET_003
+ XI1.XI0.XI1<11>.XI7<4>.NET_000 XI1.XI0.XI1<11>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_72 XI1.XI0.XI1<11>.XI7<4>.NET_007
+ XI1.XI0.XI1<11>.XI7<4>.NET_001 XI1.XI0.XI1<11>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<4>.NET_005
+ XI1.XI0.XI1<11>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<4>.NET_003
+ XI1.XI0.XI1<11>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_41_11 REG_DATA_11<11>
+ XI1.XI0.XI1<11>.XI7<11>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<11>.MM_i_7 XI1.XI0.XI1<11>.XI7<11>.NET_001
+ XI1.XI0.XI1<11>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_13 XI1.XI0.XI1<11>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_18 XI1.XI0.XI1<11>.XI7<11>.NET_003
+ XI1.XI0.XI1<11>.XI7<11>.NET_001 XI1.XI0.XI1<11>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_24 XI1.XI0.XI1<11>.XI7<11>.NET_004
+ XI1.XI0.XI1<11>.XI7<11>.NET_000 XI1.XI0.XI1<11>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<11>.NET_005
+ XI1.XI0.XI1<11>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<11>.NET_003
+ XI1.XI0.XI1<11>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_89_4 REG_DATA_11<11>
+ XI1.XI0.XI1<11>.XI7<11>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<11>.MM_i_55 XI1.XI0.XI1<11>.XI7<11>.NET_001
+ XI1.XI0.XI1<11>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_61 XI1.XI0.XI1<11>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_66 XI1.XI0.XI1<11>.XI7<11>.NET_003
+ XI1.XI0.XI1<11>.XI7<11>.NET_000 XI1.XI0.XI1<11>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_72 XI1.XI0.XI1<11>.XI7<11>.NET_007
+ XI1.XI0.XI1<11>.XI7<11>.NET_001 XI1.XI0.XI1<11>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<11>.NET_005
+ XI1.XI0.XI1<11>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<11>.NET_003
+ XI1.XI0.XI1<11>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_41_11 REG_DATA_11<10>
+ XI1.XI0.XI1<11>.XI7<10>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<10>.MM_i_7 XI1.XI0.XI1<11>.XI7<10>.NET_001
+ XI1.XI0.XI1<11>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_13 XI1.XI0.XI1<11>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_18 XI1.XI0.XI1<11>.XI7<10>.NET_003
+ XI1.XI0.XI1<11>.XI7<10>.NET_001 XI1.XI0.XI1<11>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_24 XI1.XI0.XI1<11>.XI7<10>.NET_004
+ XI1.XI0.XI1<11>.XI7<10>.NET_000 XI1.XI0.XI1<11>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<10>.NET_005
+ XI1.XI0.XI1<11>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<10>.NET_003
+ XI1.XI0.XI1<11>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_89_4 REG_DATA_11<10>
+ XI1.XI0.XI1<11>.XI7<10>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<10>.MM_i_55 XI1.XI0.XI1<11>.XI7<10>.NET_001
+ XI1.XI0.XI1<11>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_61 XI1.XI0.XI1<11>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_66 XI1.XI0.XI1<11>.XI7<10>.NET_003
+ XI1.XI0.XI1<11>.XI7<10>.NET_000 XI1.XI0.XI1<11>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_72 XI1.XI0.XI1<11>.XI7<10>.NET_007
+ XI1.XI0.XI1<11>.XI7<10>.NET_001 XI1.XI0.XI1<11>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<10>.NET_005
+ XI1.XI0.XI1<11>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<10>.NET_003
+ XI1.XI0.XI1<11>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_41_11 REG_DATA_11<9> XI1.XI0.XI1<11>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<9>.MM_i_7 XI1.XI0.XI1<11>.XI7<9>.NET_001
+ XI1.XI0.XI1<11>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_13 XI1.XI0.XI1<11>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_18 XI1.XI0.XI1<11>.XI7<9>.NET_003
+ XI1.XI0.XI1<11>.XI7<9>.NET_001 XI1.XI0.XI1<11>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_24 XI1.XI0.XI1<11>.XI7<9>.NET_004
+ XI1.XI0.XI1<11>.XI7<9>.NET_000 XI1.XI0.XI1<11>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<9>.NET_005
+ XI1.XI0.XI1<11>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<9>.NET_003
+ XI1.XI0.XI1<11>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_89_4 REG_DATA_11<9> XI1.XI0.XI1<11>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<9>.MM_i_55 XI1.XI0.XI1<11>.XI7<9>.NET_001
+ XI1.XI0.XI1<11>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_61 XI1.XI0.XI1<11>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_66 XI1.XI0.XI1<11>.XI7<9>.NET_003
+ XI1.XI0.XI1<11>.XI7<9>.NET_000 XI1.XI0.XI1<11>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_72 XI1.XI0.XI1<11>.XI7<9>.NET_007
+ XI1.XI0.XI1<11>.XI7<9>.NET_001 XI1.XI0.XI1<11>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<9>.NET_005
+ XI1.XI0.XI1<11>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<9>.NET_003
+ XI1.XI0.XI1<11>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_41_11 REG_DATA_11<8> XI1.XI0.XI1<11>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<8>.MM_i_7 XI1.XI0.XI1<11>.XI7<8>.NET_001
+ XI1.XI0.XI1<11>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_13 XI1.XI0.XI1<11>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_18 XI1.XI0.XI1<11>.XI7<8>.NET_003
+ XI1.XI0.XI1<11>.XI7<8>.NET_001 XI1.XI0.XI1<11>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_24 XI1.XI0.XI1<11>.XI7<8>.NET_004
+ XI1.XI0.XI1<11>.XI7<8>.NET_000 XI1.XI0.XI1<11>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<8>.NET_005
+ XI1.XI0.XI1<11>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<8>.NET_003
+ XI1.XI0.XI1<11>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_89_4 REG_DATA_11<8> XI1.XI0.XI1<11>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<8>.MM_i_55 XI1.XI0.XI1<11>.XI7<8>.NET_001
+ XI1.XI0.XI1<11>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_61 XI1.XI0.XI1<11>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_66 XI1.XI0.XI1<11>.XI7<8>.NET_003
+ XI1.XI0.XI1<11>.XI7<8>.NET_000 XI1.XI0.XI1<11>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_72 XI1.XI0.XI1<11>.XI7<8>.NET_007
+ XI1.XI0.XI1<11>.XI7<8>.NET_001 XI1.XI0.XI1<11>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<8>.NET_005
+ XI1.XI0.XI1<11>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<8>.NET_003
+ XI1.XI0.XI1<11>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_41_11 REG_DATA_11<15>
+ XI1.XI0.XI1<11>.XI7<15>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<15>.MM_i_7 XI1.XI0.XI1<11>.XI7<15>.NET_001
+ XI1.XI0.XI1<11>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_13 XI1.XI0.XI1<11>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_18 XI1.XI0.XI1<11>.XI7<15>.NET_003
+ XI1.XI0.XI1<11>.XI7<15>.NET_001 XI1.XI0.XI1<11>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_24 XI1.XI0.XI1<11>.XI7<15>.NET_004
+ XI1.XI0.XI1<11>.XI7<15>.NET_000 XI1.XI0.XI1<11>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<15>.NET_005
+ XI1.XI0.XI1<11>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<15>.NET_003
+ XI1.XI0.XI1<11>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_89_4 REG_DATA_11<15>
+ XI1.XI0.XI1<11>.XI7<15>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<15>.MM_i_55 XI1.XI0.XI1<11>.XI7<15>.NET_001
+ XI1.XI0.XI1<11>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_61 XI1.XI0.XI1<11>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_66 XI1.XI0.XI1<11>.XI7<15>.NET_003
+ XI1.XI0.XI1<11>.XI7<15>.NET_000 XI1.XI0.XI1<11>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_72 XI1.XI0.XI1<11>.XI7<15>.NET_007
+ XI1.XI0.XI1<11>.XI7<15>.NET_001 XI1.XI0.XI1<11>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<15>.NET_005
+ XI1.XI0.XI1<11>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<15>.NET_003
+ XI1.XI0.XI1<11>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_41_11 REG_DATA_11<14>
+ XI1.XI0.XI1<11>.XI7<14>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<14>.MM_i_7 XI1.XI0.XI1<11>.XI7<14>.NET_001
+ XI1.XI0.XI1<11>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_13 XI1.XI0.XI1<11>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_18 XI1.XI0.XI1<11>.XI7<14>.NET_003
+ XI1.XI0.XI1<11>.XI7<14>.NET_001 XI1.XI0.XI1<11>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_24 XI1.XI0.XI1<11>.XI7<14>.NET_004
+ XI1.XI0.XI1<11>.XI7<14>.NET_000 XI1.XI0.XI1<11>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<14>.NET_005
+ XI1.XI0.XI1<11>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<14>.NET_003
+ XI1.XI0.XI1<11>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_89_4 REG_DATA_11<14>
+ XI1.XI0.XI1<11>.XI7<14>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<14>.MM_i_55 XI1.XI0.XI1<11>.XI7<14>.NET_001
+ XI1.XI0.XI1<11>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_61 XI1.XI0.XI1<11>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_66 XI1.XI0.XI1<11>.XI7<14>.NET_003
+ XI1.XI0.XI1<11>.XI7<14>.NET_000 XI1.XI0.XI1<11>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_72 XI1.XI0.XI1<11>.XI7<14>.NET_007
+ XI1.XI0.XI1<11>.XI7<14>.NET_001 XI1.XI0.XI1<11>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<14>.NET_005
+ XI1.XI0.XI1<11>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<14>.NET_003
+ XI1.XI0.XI1<11>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_41_11 REG_DATA_11<13>
+ XI1.XI0.XI1<11>.XI7<13>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<13>.MM_i_7 XI1.XI0.XI1<11>.XI7<13>.NET_001
+ XI1.XI0.XI1<11>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_13 XI1.XI0.XI1<11>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_18 XI1.XI0.XI1<11>.XI7<13>.NET_003
+ XI1.XI0.XI1<11>.XI7<13>.NET_001 XI1.XI0.XI1<11>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_24 XI1.XI0.XI1<11>.XI7<13>.NET_004
+ XI1.XI0.XI1<11>.XI7<13>.NET_000 XI1.XI0.XI1<11>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<13>.NET_005
+ XI1.XI0.XI1<11>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<13>.NET_003
+ XI1.XI0.XI1<11>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_89_4 REG_DATA_11<13>
+ XI1.XI0.XI1<11>.XI7<13>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<13>.MM_i_55 XI1.XI0.XI1<11>.XI7<13>.NET_001
+ XI1.XI0.XI1<11>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_61 XI1.XI0.XI1<11>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_66 XI1.XI0.XI1<11>.XI7<13>.NET_003
+ XI1.XI0.XI1<11>.XI7<13>.NET_000 XI1.XI0.XI1<11>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_72 XI1.XI0.XI1<11>.XI7<13>.NET_007
+ XI1.XI0.XI1<11>.XI7<13>.NET_001 XI1.XI0.XI1<11>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<13>.NET_005
+ XI1.XI0.XI1<11>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<13>.NET_003
+ XI1.XI0.XI1<11>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_41_11 REG_DATA_11<12>
+ XI1.XI0.XI1<11>.XI7<12>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<11>.XI7<12>.MM_i_7 XI1.XI0.XI1<11>.XI7<12>.NET_001
+ XI1.XI0.XI1<11>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_13 XI1.XI0.XI1<11>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_18 XI1.XI0.XI1<11>.XI7<12>.NET_003
+ XI1.XI0.XI1<11>.XI7<12>.NET_001 XI1.XI0.XI1<11>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_24 XI1.XI0.XI1<11>.XI7<12>.NET_004
+ XI1.XI0.XI1<11>.XI7<12>.NET_000 XI1.XI0.XI1<11>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<11>.XI7<12>.NET_005
+ XI1.XI0.XI1<11>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<11>.XI7<12>.NET_003
+ XI1.XI0.XI1<11>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<11>
+ XI1.XI0.XI1<11>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_89_4 REG_DATA_11<12>
+ XI1.XI0.XI1<11>.XI7<12>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<11>.XI7<12>.MM_i_55 XI1.XI0.XI1<11>.XI7<12>.NET_001
+ XI1.XI0.XI1<11>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_61 XI1.XI0.XI1<11>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_66 XI1.XI0.XI1<11>.XI7<12>.NET_003
+ XI1.XI0.XI1<11>.XI7<12>.NET_000 XI1.XI0.XI1<11>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_72 XI1.XI0.XI1<11>.XI7<12>.NET_007
+ XI1.XI0.XI1<11>.XI7<12>.NET_001 XI1.XI0.XI1<11>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<11>.XI7<12>.NET_005
+ XI1.XI0.XI1<11>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<11>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<11>.XI7<12>.NET_003
+ XI1.XI0.XI1<11>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_41_11 REG_DATA_10<3> XI1.XI0.XI1<10>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<3>.MM_i_7 XI1.XI0.XI1<10>.XI7<3>.NET_001
+ XI1.XI0.XI1<10>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_13 XI1.XI0.XI1<10>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_18 XI1.XI0.XI1<10>.XI7<3>.NET_003
+ XI1.XI0.XI1<10>.XI7<3>.NET_001 XI1.XI0.XI1<10>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_24 XI1.XI0.XI1<10>.XI7<3>.NET_004
+ XI1.XI0.XI1<10>.XI7<3>.NET_000 XI1.XI0.XI1<10>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<3>.NET_005
+ XI1.XI0.XI1<10>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<3>.NET_003
+ XI1.XI0.XI1<10>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_89_4 REG_DATA_10<3> XI1.XI0.XI1<10>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<3>.MM_i_55 XI1.XI0.XI1<10>.XI7<3>.NET_001
+ XI1.XI0.XI1<10>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_61 XI1.XI0.XI1<10>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_66 XI1.XI0.XI1<10>.XI7<3>.NET_003
+ XI1.XI0.XI1<10>.XI7<3>.NET_000 XI1.XI0.XI1<10>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_72 XI1.XI0.XI1<10>.XI7<3>.NET_007
+ XI1.XI0.XI1<10>.XI7<3>.NET_001 XI1.XI0.XI1<10>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<3>.NET_005
+ XI1.XI0.XI1<10>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<3>.NET_003
+ XI1.XI0.XI1<10>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_41_11 REG_DATA_10<2> XI1.XI0.XI1<10>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<2>.MM_i_7 XI1.XI0.XI1<10>.XI7<2>.NET_001
+ XI1.XI0.XI1<10>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_13 XI1.XI0.XI1<10>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_18 XI1.XI0.XI1<10>.XI7<2>.NET_003
+ XI1.XI0.XI1<10>.XI7<2>.NET_001 XI1.XI0.XI1<10>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_24 XI1.XI0.XI1<10>.XI7<2>.NET_004
+ XI1.XI0.XI1<10>.XI7<2>.NET_000 XI1.XI0.XI1<10>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<2>.NET_005
+ XI1.XI0.XI1<10>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<2>.NET_003
+ XI1.XI0.XI1<10>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_89_4 REG_DATA_10<2> XI1.XI0.XI1<10>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<2>.MM_i_55 XI1.XI0.XI1<10>.XI7<2>.NET_001
+ XI1.XI0.XI1<10>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_61 XI1.XI0.XI1<10>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_66 XI1.XI0.XI1<10>.XI7<2>.NET_003
+ XI1.XI0.XI1<10>.XI7<2>.NET_000 XI1.XI0.XI1<10>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_72 XI1.XI0.XI1<10>.XI7<2>.NET_007
+ XI1.XI0.XI1<10>.XI7<2>.NET_001 XI1.XI0.XI1<10>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<2>.NET_005
+ XI1.XI0.XI1<10>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<2>.NET_003
+ XI1.XI0.XI1<10>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_41_11 REG_DATA_10<1> XI1.XI0.XI1<10>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<1>.MM_i_7 XI1.XI0.XI1<10>.XI7<1>.NET_001
+ XI1.XI0.XI1<10>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_13 XI1.XI0.XI1<10>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_18 XI1.XI0.XI1<10>.XI7<1>.NET_003
+ XI1.XI0.XI1<10>.XI7<1>.NET_001 XI1.XI0.XI1<10>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_24 XI1.XI0.XI1<10>.XI7<1>.NET_004
+ XI1.XI0.XI1<10>.XI7<1>.NET_000 XI1.XI0.XI1<10>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<1>.NET_005
+ XI1.XI0.XI1<10>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<1>.NET_003
+ XI1.XI0.XI1<10>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_89_4 REG_DATA_10<1> XI1.XI0.XI1<10>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<1>.MM_i_55 XI1.XI0.XI1<10>.XI7<1>.NET_001
+ XI1.XI0.XI1<10>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_61 XI1.XI0.XI1<10>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_66 XI1.XI0.XI1<10>.XI7<1>.NET_003
+ XI1.XI0.XI1<10>.XI7<1>.NET_000 XI1.XI0.XI1<10>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_72 XI1.XI0.XI1<10>.XI7<1>.NET_007
+ XI1.XI0.XI1<10>.XI7<1>.NET_001 XI1.XI0.XI1<10>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<1>.NET_005
+ XI1.XI0.XI1<10>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<1>.NET_003
+ XI1.XI0.XI1<10>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_41_11 REG_DATA_10<0> XI1.XI0.XI1<10>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<0>.MM_i_7 XI1.XI0.XI1<10>.XI7<0>.NET_001
+ XI1.XI0.XI1<10>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_13 XI1.XI0.XI1<10>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_18 XI1.XI0.XI1<10>.XI7<0>.NET_003
+ XI1.XI0.XI1<10>.XI7<0>.NET_001 XI1.XI0.XI1<10>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_24 XI1.XI0.XI1<10>.XI7<0>.NET_004
+ XI1.XI0.XI1<10>.XI7<0>.NET_000 XI1.XI0.XI1<10>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<0>.NET_005
+ XI1.XI0.XI1<10>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<0>.NET_003
+ XI1.XI0.XI1<10>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_89_4 REG_DATA_10<0> XI1.XI0.XI1<10>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<0>.MM_i_55 XI1.XI0.XI1<10>.XI7<0>.NET_001
+ XI1.XI0.XI1<10>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_61 XI1.XI0.XI1<10>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_66 XI1.XI0.XI1<10>.XI7<0>.NET_003
+ XI1.XI0.XI1<10>.XI7<0>.NET_000 XI1.XI0.XI1<10>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_72 XI1.XI0.XI1<10>.XI7<0>.NET_007
+ XI1.XI0.XI1<10>.XI7<0>.NET_001 XI1.XI0.XI1<10>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<0>.NET_005
+ XI1.XI0.XI1<10>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<0>.NET_003
+ XI1.XI0.XI1<10>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_41_11 REG_DATA_10<7> XI1.XI0.XI1<10>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<7>.MM_i_7 XI1.XI0.XI1<10>.XI7<7>.NET_001
+ XI1.XI0.XI1<10>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_13 XI1.XI0.XI1<10>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_18 XI1.XI0.XI1<10>.XI7<7>.NET_003
+ XI1.XI0.XI1<10>.XI7<7>.NET_001 XI1.XI0.XI1<10>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_24 XI1.XI0.XI1<10>.XI7<7>.NET_004
+ XI1.XI0.XI1<10>.XI7<7>.NET_000 XI1.XI0.XI1<10>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<7>.NET_005
+ XI1.XI0.XI1<10>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<7>.NET_003
+ XI1.XI0.XI1<10>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_89_4 REG_DATA_10<7> XI1.XI0.XI1<10>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<7>.MM_i_55 XI1.XI0.XI1<10>.XI7<7>.NET_001
+ XI1.XI0.XI1<10>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_61 XI1.XI0.XI1<10>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_66 XI1.XI0.XI1<10>.XI7<7>.NET_003
+ XI1.XI0.XI1<10>.XI7<7>.NET_000 XI1.XI0.XI1<10>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_72 XI1.XI0.XI1<10>.XI7<7>.NET_007
+ XI1.XI0.XI1<10>.XI7<7>.NET_001 XI1.XI0.XI1<10>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<7>.NET_005
+ XI1.XI0.XI1<10>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<7>.NET_003
+ XI1.XI0.XI1<10>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_41_11 REG_DATA_10<6> XI1.XI0.XI1<10>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<6>.MM_i_7 XI1.XI0.XI1<10>.XI7<6>.NET_001
+ XI1.XI0.XI1<10>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_13 XI1.XI0.XI1<10>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_18 XI1.XI0.XI1<10>.XI7<6>.NET_003
+ XI1.XI0.XI1<10>.XI7<6>.NET_001 XI1.XI0.XI1<10>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_24 XI1.XI0.XI1<10>.XI7<6>.NET_004
+ XI1.XI0.XI1<10>.XI7<6>.NET_000 XI1.XI0.XI1<10>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<6>.NET_005
+ XI1.XI0.XI1<10>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<6>.NET_003
+ XI1.XI0.XI1<10>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_89_4 REG_DATA_10<6> XI1.XI0.XI1<10>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<6>.MM_i_55 XI1.XI0.XI1<10>.XI7<6>.NET_001
+ XI1.XI0.XI1<10>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_61 XI1.XI0.XI1<10>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_66 XI1.XI0.XI1<10>.XI7<6>.NET_003
+ XI1.XI0.XI1<10>.XI7<6>.NET_000 XI1.XI0.XI1<10>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_72 XI1.XI0.XI1<10>.XI7<6>.NET_007
+ XI1.XI0.XI1<10>.XI7<6>.NET_001 XI1.XI0.XI1<10>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<6>.NET_005
+ XI1.XI0.XI1<10>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<6>.NET_003
+ XI1.XI0.XI1<10>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_41_11 REG_DATA_10<5> XI1.XI0.XI1<10>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<5>.MM_i_7 XI1.XI0.XI1<10>.XI7<5>.NET_001
+ XI1.XI0.XI1<10>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_13 XI1.XI0.XI1<10>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_18 XI1.XI0.XI1<10>.XI7<5>.NET_003
+ XI1.XI0.XI1<10>.XI7<5>.NET_001 XI1.XI0.XI1<10>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_24 XI1.XI0.XI1<10>.XI7<5>.NET_004
+ XI1.XI0.XI1<10>.XI7<5>.NET_000 XI1.XI0.XI1<10>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<5>.NET_005
+ XI1.XI0.XI1<10>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<5>.NET_003
+ XI1.XI0.XI1<10>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_89_4 REG_DATA_10<5> XI1.XI0.XI1<10>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<5>.MM_i_55 XI1.XI0.XI1<10>.XI7<5>.NET_001
+ XI1.XI0.XI1<10>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_61 XI1.XI0.XI1<10>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_66 XI1.XI0.XI1<10>.XI7<5>.NET_003
+ XI1.XI0.XI1<10>.XI7<5>.NET_000 XI1.XI0.XI1<10>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_72 XI1.XI0.XI1<10>.XI7<5>.NET_007
+ XI1.XI0.XI1<10>.XI7<5>.NET_001 XI1.XI0.XI1<10>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<5>.NET_005
+ XI1.XI0.XI1<10>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<5>.NET_003
+ XI1.XI0.XI1<10>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_41_11 REG_DATA_10<4> XI1.XI0.XI1<10>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<4>.MM_i_7 XI1.XI0.XI1<10>.XI7<4>.NET_001
+ XI1.XI0.XI1<10>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_13 XI1.XI0.XI1<10>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_18 XI1.XI0.XI1<10>.XI7<4>.NET_003
+ XI1.XI0.XI1<10>.XI7<4>.NET_001 XI1.XI0.XI1<10>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_24 XI1.XI0.XI1<10>.XI7<4>.NET_004
+ XI1.XI0.XI1<10>.XI7<4>.NET_000 XI1.XI0.XI1<10>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<4>.NET_005
+ XI1.XI0.XI1<10>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<4>.NET_003
+ XI1.XI0.XI1<10>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_89_4 REG_DATA_10<4> XI1.XI0.XI1<10>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<4>.MM_i_55 XI1.XI0.XI1<10>.XI7<4>.NET_001
+ XI1.XI0.XI1<10>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_61 XI1.XI0.XI1<10>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_66 XI1.XI0.XI1<10>.XI7<4>.NET_003
+ XI1.XI0.XI1<10>.XI7<4>.NET_000 XI1.XI0.XI1<10>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_72 XI1.XI0.XI1<10>.XI7<4>.NET_007
+ XI1.XI0.XI1<10>.XI7<4>.NET_001 XI1.XI0.XI1<10>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<4>.NET_005
+ XI1.XI0.XI1<10>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<4>.NET_003
+ XI1.XI0.XI1<10>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_41_11 REG_DATA_10<11>
+ XI1.XI0.XI1<10>.XI7<11>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<11>.MM_i_7 XI1.XI0.XI1<10>.XI7<11>.NET_001
+ XI1.XI0.XI1<10>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_13 XI1.XI0.XI1<10>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_18 XI1.XI0.XI1<10>.XI7<11>.NET_003
+ XI1.XI0.XI1<10>.XI7<11>.NET_001 XI1.XI0.XI1<10>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_24 XI1.XI0.XI1<10>.XI7<11>.NET_004
+ XI1.XI0.XI1<10>.XI7<11>.NET_000 XI1.XI0.XI1<10>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<11>.NET_005
+ XI1.XI0.XI1<10>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<11>.NET_003
+ XI1.XI0.XI1<10>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_89_4 REG_DATA_10<11>
+ XI1.XI0.XI1<10>.XI7<11>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<11>.MM_i_55 XI1.XI0.XI1<10>.XI7<11>.NET_001
+ XI1.XI0.XI1<10>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_61 XI1.XI0.XI1<10>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_66 XI1.XI0.XI1<10>.XI7<11>.NET_003
+ XI1.XI0.XI1<10>.XI7<11>.NET_000 XI1.XI0.XI1<10>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_72 XI1.XI0.XI1<10>.XI7<11>.NET_007
+ XI1.XI0.XI1<10>.XI7<11>.NET_001 XI1.XI0.XI1<10>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<11>.NET_005
+ XI1.XI0.XI1<10>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<11>.NET_003
+ XI1.XI0.XI1<10>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_41_11 REG_DATA_10<10>
+ XI1.XI0.XI1<10>.XI7<10>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<10>.MM_i_7 XI1.XI0.XI1<10>.XI7<10>.NET_001
+ XI1.XI0.XI1<10>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_13 XI1.XI0.XI1<10>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_18 XI1.XI0.XI1<10>.XI7<10>.NET_003
+ XI1.XI0.XI1<10>.XI7<10>.NET_001 XI1.XI0.XI1<10>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_24 XI1.XI0.XI1<10>.XI7<10>.NET_004
+ XI1.XI0.XI1<10>.XI7<10>.NET_000 XI1.XI0.XI1<10>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<10>.NET_005
+ XI1.XI0.XI1<10>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<10>.NET_003
+ XI1.XI0.XI1<10>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_89_4 REG_DATA_10<10>
+ XI1.XI0.XI1<10>.XI7<10>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<10>.MM_i_55 XI1.XI0.XI1<10>.XI7<10>.NET_001
+ XI1.XI0.XI1<10>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_61 XI1.XI0.XI1<10>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_66 XI1.XI0.XI1<10>.XI7<10>.NET_003
+ XI1.XI0.XI1<10>.XI7<10>.NET_000 XI1.XI0.XI1<10>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_72 XI1.XI0.XI1<10>.XI7<10>.NET_007
+ XI1.XI0.XI1<10>.XI7<10>.NET_001 XI1.XI0.XI1<10>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<10>.NET_005
+ XI1.XI0.XI1<10>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<10>.NET_003
+ XI1.XI0.XI1<10>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_41_11 REG_DATA_10<9> XI1.XI0.XI1<10>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<9>.MM_i_7 XI1.XI0.XI1<10>.XI7<9>.NET_001
+ XI1.XI0.XI1<10>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_13 XI1.XI0.XI1<10>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_18 XI1.XI0.XI1<10>.XI7<9>.NET_003
+ XI1.XI0.XI1<10>.XI7<9>.NET_001 XI1.XI0.XI1<10>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_24 XI1.XI0.XI1<10>.XI7<9>.NET_004
+ XI1.XI0.XI1<10>.XI7<9>.NET_000 XI1.XI0.XI1<10>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<9>.NET_005
+ XI1.XI0.XI1<10>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<9>.NET_003
+ XI1.XI0.XI1<10>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_89_4 REG_DATA_10<9> XI1.XI0.XI1<10>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<9>.MM_i_55 XI1.XI0.XI1<10>.XI7<9>.NET_001
+ XI1.XI0.XI1<10>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_61 XI1.XI0.XI1<10>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_66 XI1.XI0.XI1<10>.XI7<9>.NET_003
+ XI1.XI0.XI1<10>.XI7<9>.NET_000 XI1.XI0.XI1<10>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_72 XI1.XI0.XI1<10>.XI7<9>.NET_007
+ XI1.XI0.XI1<10>.XI7<9>.NET_001 XI1.XI0.XI1<10>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<9>.NET_005
+ XI1.XI0.XI1<10>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<9>.NET_003
+ XI1.XI0.XI1<10>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_41_11 REG_DATA_10<8> XI1.XI0.XI1<10>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<8>.MM_i_7 XI1.XI0.XI1<10>.XI7<8>.NET_001
+ XI1.XI0.XI1<10>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_13 XI1.XI0.XI1<10>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_18 XI1.XI0.XI1<10>.XI7<8>.NET_003
+ XI1.XI0.XI1<10>.XI7<8>.NET_001 XI1.XI0.XI1<10>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_24 XI1.XI0.XI1<10>.XI7<8>.NET_004
+ XI1.XI0.XI1<10>.XI7<8>.NET_000 XI1.XI0.XI1<10>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<8>.NET_005
+ XI1.XI0.XI1<10>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<8>.NET_003
+ XI1.XI0.XI1<10>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_89_4 REG_DATA_10<8> XI1.XI0.XI1<10>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<8>.MM_i_55 XI1.XI0.XI1<10>.XI7<8>.NET_001
+ XI1.XI0.XI1<10>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_61 XI1.XI0.XI1<10>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_66 XI1.XI0.XI1<10>.XI7<8>.NET_003
+ XI1.XI0.XI1<10>.XI7<8>.NET_000 XI1.XI0.XI1<10>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_72 XI1.XI0.XI1<10>.XI7<8>.NET_007
+ XI1.XI0.XI1<10>.XI7<8>.NET_001 XI1.XI0.XI1<10>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<8>.NET_005
+ XI1.XI0.XI1<10>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<8>.NET_003
+ XI1.XI0.XI1<10>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_41_11 REG_DATA_10<15>
+ XI1.XI0.XI1<10>.XI7<15>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<15>.MM_i_7 XI1.XI0.XI1<10>.XI7<15>.NET_001
+ XI1.XI0.XI1<10>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_13 XI1.XI0.XI1<10>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_18 XI1.XI0.XI1<10>.XI7<15>.NET_003
+ XI1.XI0.XI1<10>.XI7<15>.NET_001 XI1.XI0.XI1<10>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_24 XI1.XI0.XI1<10>.XI7<15>.NET_004
+ XI1.XI0.XI1<10>.XI7<15>.NET_000 XI1.XI0.XI1<10>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<15>.NET_005
+ XI1.XI0.XI1<10>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<15>.NET_003
+ XI1.XI0.XI1<10>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_89_4 REG_DATA_10<15>
+ XI1.XI0.XI1<10>.XI7<15>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<15>.MM_i_55 XI1.XI0.XI1<10>.XI7<15>.NET_001
+ XI1.XI0.XI1<10>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_61 XI1.XI0.XI1<10>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_66 XI1.XI0.XI1<10>.XI7<15>.NET_003
+ XI1.XI0.XI1<10>.XI7<15>.NET_000 XI1.XI0.XI1<10>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_72 XI1.XI0.XI1<10>.XI7<15>.NET_007
+ XI1.XI0.XI1<10>.XI7<15>.NET_001 XI1.XI0.XI1<10>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<15>.NET_005
+ XI1.XI0.XI1<10>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<15>.NET_003
+ XI1.XI0.XI1<10>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_41_11 REG_DATA_10<14>
+ XI1.XI0.XI1<10>.XI7<14>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<14>.MM_i_7 XI1.XI0.XI1<10>.XI7<14>.NET_001
+ XI1.XI0.XI1<10>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_13 XI1.XI0.XI1<10>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_18 XI1.XI0.XI1<10>.XI7<14>.NET_003
+ XI1.XI0.XI1<10>.XI7<14>.NET_001 XI1.XI0.XI1<10>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_24 XI1.XI0.XI1<10>.XI7<14>.NET_004
+ XI1.XI0.XI1<10>.XI7<14>.NET_000 XI1.XI0.XI1<10>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<14>.NET_005
+ XI1.XI0.XI1<10>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<14>.NET_003
+ XI1.XI0.XI1<10>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_89_4 REG_DATA_10<14>
+ XI1.XI0.XI1<10>.XI7<14>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<14>.MM_i_55 XI1.XI0.XI1<10>.XI7<14>.NET_001
+ XI1.XI0.XI1<10>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_61 XI1.XI0.XI1<10>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_66 XI1.XI0.XI1<10>.XI7<14>.NET_003
+ XI1.XI0.XI1<10>.XI7<14>.NET_000 XI1.XI0.XI1<10>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_72 XI1.XI0.XI1<10>.XI7<14>.NET_007
+ XI1.XI0.XI1<10>.XI7<14>.NET_001 XI1.XI0.XI1<10>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<14>.NET_005
+ XI1.XI0.XI1<10>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<14>.NET_003
+ XI1.XI0.XI1<10>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_41_11 REG_DATA_10<13>
+ XI1.XI0.XI1<10>.XI7<13>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<13>.MM_i_7 XI1.XI0.XI1<10>.XI7<13>.NET_001
+ XI1.XI0.XI1<10>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_13 XI1.XI0.XI1<10>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_18 XI1.XI0.XI1<10>.XI7<13>.NET_003
+ XI1.XI0.XI1<10>.XI7<13>.NET_001 XI1.XI0.XI1<10>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_24 XI1.XI0.XI1<10>.XI7<13>.NET_004
+ XI1.XI0.XI1<10>.XI7<13>.NET_000 XI1.XI0.XI1<10>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<13>.NET_005
+ XI1.XI0.XI1<10>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<13>.NET_003
+ XI1.XI0.XI1<10>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_89_4 REG_DATA_10<13>
+ XI1.XI0.XI1<10>.XI7<13>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<13>.MM_i_55 XI1.XI0.XI1<10>.XI7<13>.NET_001
+ XI1.XI0.XI1<10>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_61 XI1.XI0.XI1<10>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_66 XI1.XI0.XI1<10>.XI7<13>.NET_003
+ XI1.XI0.XI1<10>.XI7<13>.NET_000 XI1.XI0.XI1<10>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_72 XI1.XI0.XI1<10>.XI7<13>.NET_007
+ XI1.XI0.XI1<10>.XI7<13>.NET_001 XI1.XI0.XI1<10>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<13>.NET_005
+ XI1.XI0.XI1<10>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<13>.NET_003
+ XI1.XI0.XI1<10>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_41_11 REG_DATA_10<12>
+ XI1.XI0.XI1<10>.XI7<12>.NET_003 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI1<10>.XI7<12>.MM_i_7 XI1.XI0.XI1<10>.XI7<12>.NET_001
+ XI1.XI0.XI1<10>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_13 XI1.XI0.XI1<10>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_18 XI1.XI0.XI1<10>.XI7<12>.NET_003
+ XI1.XI0.XI1<10>.XI7<12>.NET_001 XI1.XI0.XI1<10>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_24 XI1.XI0.XI1<10>.XI7<12>.NET_004
+ XI1.XI0.XI1<10>.XI7<12>.NET_000 XI1.XI0.XI1<10>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<10>.XI7<12>.NET_005
+ XI1.XI0.XI1<10>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<10>.XI7<12>.NET_003
+ XI1.XI0.XI1<10>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<10>
+ XI1.XI0.XI1<10>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_89_4 REG_DATA_10<12>
+ XI1.XI0.XI1<10>.XI7<12>.NET_003 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI1<10>.XI7<12>.MM_i_55 XI1.XI0.XI1<10>.XI7<12>.NET_001
+ XI1.XI0.XI1<10>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_61 XI1.XI0.XI1<10>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_66 XI1.XI0.XI1<10>.XI7<12>.NET_003
+ XI1.XI0.XI1<10>.XI7<12>.NET_000 XI1.XI0.XI1<10>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_72 XI1.XI0.XI1<10>.XI7<12>.NET_007
+ XI1.XI0.XI1<10>.XI7<12>.NET_001 XI1.XI0.XI1<10>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<10>.XI7<12>.NET_005
+ XI1.XI0.XI1<10>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<10>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<10>.XI7<12>.NET_003
+ XI1.XI0.XI1<10>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_41_11 REG_DATA_9<3> XI1.XI0.XI1<9>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<3>.MM_i_7 XI1.XI0.XI1<9>.XI7<3>.NET_001
+ XI1.XI0.XI1<9>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_13 XI1.XI0.XI1<9>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_18 XI1.XI0.XI1<9>.XI7<3>.NET_003
+ XI1.XI0.XI1<9>.XI7<3>.NET_001 XI1.XI0.XI1<9>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_24 XI1.XI0.XI1<9>.XI7<3>.NET_004
+ XI1.XI0.XI1<9>.XI7<3>.NET_000 XI1.XI0.XI1<9>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<3>.NET_005
+ XI1.XI0.XI1<9>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<3>.NET_003
+ XI1.XI0.XI1<9>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_89_4 REG_DATA_9<3> XI1.XI0.XI1<9>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<3>.MM_i_55 XI1.XI0.XI1<9>.XI7<3>.NET_001
+ XI1.XI0.XI1<9>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_61 XI1.XI0.XI1<9>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_66 XI1.XI0.XI1<9>.XI7<3>.NET_003
+ XI1.XI0.XI1<9>.XI7<3>.NET_000 XI1.XI0.XI1<9>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_72 XI1.XI0.XI1<9>.XI7<3>.NET_007
+ XI1.XI0.XI1<9>.XI7<3>.NET_001 XI1.XI0.XI1<9>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<3>.NET_005
+ XI1.XI0.XI1<9>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<3>.NET_003
+ XI1.XI0.XI1<9>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_41_11 REG_DATA_9<2> XI1.XI0.XI1<9>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<2>.MM_i_7 XI1.XI0.XI1<9>.XI7<2>.NET_001
+ XI1.XI0.XI1<9>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_13 XI1.XI0.XI1<9>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_18 XI1.XI0.XI1<9>.XI7<2>.NET_003
+ XI1.XI0.XI1<9>.XI7<2>.NET_001 XI1.XI0.XI1<9>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_24 XI1.XI0.XI1<9>.XI7<2>.NET_004
+ XI1.XI0.XI1<9>.XI7<2>.NET_000 XI1.XI0.XI1<9>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<2>.NET_005
+ XI1.XI0.XI1<9>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<2>.NET_003
+ XI1.XI0.XI1<9>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_89_4 REG_DATA_9<2> XI1.XI0.XI1<9>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<2>.MM_i_55 XI1.XI0.XI1<9>.XI7<2>.NET_001
+ XI1.XI0.XI1<9>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_61 XI1.XI0.XI1<9>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_66 XI1.XI0.XI1<9>.XI7<2>.NET_003
+ XI1.XI0.XI1<9>.XI7<2>.NET_000 XI1.XI0.XI1<9>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_72 XI1.XI0.XI1<9>.XI7<2>.NET_007
+ XI1.XI0.XI1<9>.XI7<2>.NET_001 XI1.XI0.XI1<9>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<2>.NET_005
+ XI1.XI0.XI1<9>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<2>.NET_003
+ XI1.XI0.XI1<9>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_41_11 REG_DATA_9<1> XI1.XI0.XI1<9>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<1>.MM_i_7 XI1.XI0.XI1<9>.XI7<1>.NET_001
+ XI1.XI0.XI1<9>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_13 XI1.XI0.XI1<9>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_18 XI1.XI0.XI1<9>.XI7<1>.NET_003
+ XI1.XI0.XI1<9>.XI7<1>.NET_001 XI1.XI0.XI1<9>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_24 XI1.XI0.XI1<9>.XI7<1>.NET_004
+ XI1.XI0.XI1<9>.XI7<1>.NET_000 XI1.XI0.XI1<9>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<1>.NET_005
+ XI1.XI0.XI1<9>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<1>.NET_003
+ XI1.XI0.XI1<9>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_89_4 REG_DATA_9<1> XI1.XI0.XI1<9>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<1>.MM_i_55 XI1.XI0.XI1<9>.XI7<1>.NET_001
+ XI1.XI0.XI1<9>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_61 XI1.XI0.XI1<9>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_66 XI1.XI0.XI1<9>.XI7<1>.NET_003
+ XI1.XI0.XI1<9>.XI7<1>.NET_000 XI1.XI0.XI1<9>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_72 XI1.XI0.XI1<9>.XI7<1>.NET_007
+ XI1.XI0.XI1<9>.XI7<1>.NET_001 XI1.XI0.XI1<9>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<1>.NET_005
+ XI1.XI0.XI1<9>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<1>.NET_003
+ XI1.XI0.XI1<9>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_41_11 REG_DATA_9<0> XI1.XI0.XI1<9>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<0>.MM_i_7 XI1.XI0.XI1<9>.XI7<0>.NET_001
+ XI1.XI0.XI1<9>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_13 XI1.XI0.XI1<9>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_18 XI1.XI0.XI1<9>.XI7<0>.NET_003
+ XI1.XI0.XI1<9>.XI7<0>.NET_001 XI1.XI0.XI1<9>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_24 XI1.XI0.XI1<9>.XI7<0>.NET_004
+ XI1.XI0.XI1<9>.XI7<0>.NET_000 XI1.XI0.XI1<9>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<0>.NET_005
+ XI1.XI0.XI1<9>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<0>.NET_003
+ XI1.XI0.XI1<9>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_89_4 REG_DATA_9<0> XI1.XI0.XI1<9>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<0>.MM_i_55 XI1.XI0.XI1<9>.XI7<0>.NET_001
+ XI1.XI0.XI1<9>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_61 XI1.XI0.XI1<9>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_66 XI1.XI0.XI1<9>.XI7<0>.NET_003
+ XI1.XI0.XI1<9>.XI7<0>.NET_000 XI1.XI0.XI1<9>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_72 XI1.XI0.XI1<9>.XI7<0>.NET_007
+ XI1.XI0.XI1<9>.XI7<0>.NET_001 XI1.XI0.XI1<9>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<0>.NET_005
+ XI1.XI0.XI1<9>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<0>.NET_003
+ XI1.XI0.XI1<9>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_41_11 REG_DATA_9<7> XI1.XI0.XI1<9>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<7>.MM_i_7 XI1.XI0.XI1<9>.XI7<7>.NET_001
+ XI1.XI0.XI1<9>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_13 XI1.XI0.XI1<9>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_18 XI1.XI0.XI1<9>.XI7<7>.NET_003
+ XI1.XI0.XI1<9>.XI7<7>.NET_001 XI1.XI0.XI1<9>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_24 XI1.XI0.XI1<9>.XI7<7>.NET_004
+ XI1.XI0.XI1<9>.XI7<7>.NET_000 XI1.XI0.XI1<9>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<7>.NET_005
+ XI1.XI0.XI1<9>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<7>.NET_003
+ XI1.XI0.XI1<9>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_89_4 REG_DATA_9<7> XI1.XI0.XI1<9>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<7>.MM_i_55 XI1.XI0.XI1<9>.XI7<7>.NET_001
+ XI1.XI0.XI1<9>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_61 XI1.XI0.XI1<9>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_66 XI1.XI0.XI1<9>.XI7<7>.NET_003
+ XI1.XI0.XI1<9>.XI7<7>.NET_000 XI1.XI0.XI1<9>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_72 XI1.XI0.XI1<9>.XI7<7>.NET_007
+ XI1.XI0.XI1<9>.XI7<7>.NET_001 XI1.XI0.XI1<9>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<7>.NET_005
+ XI1.XI0.XI1<9>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<7>.NET_003
+ XI1.XI0.XI1<9>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_41_11 REG_DATA_9<6> XI1.XI0.XI1<9>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<6>.MM_i_7 XI1.XI0.XI1<9>.XI7<6>.NET_001
+ XI1.XI0.XI1<9>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_13 XI1.XI0.XI1<9>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_18 XI1.XI0.XI1<9>.XI7<6>.NET_003
+ XI1.XI0.XI1<9>.XI7<6>.NET_001 XI1.XI0.XI1<9>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_24 XI1.XI0.XI1<9>.XI7<6>.NET_004
+ XI1.XI0.XI1<9>.XI7<6>.NET_000 XI1.XI0.XI1<9>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<6>.NET_005
+ XI1.XI0.XI1<9>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<6>.NET_003
+ XI1.XI0.XI1<9>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_89_4 REG_DATA_9<6> XI1.XI0.XI1<9>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<6>.MM_i_55 XI1.XI0.XI1<9>.XI7<6>.NET_001
+ XI1.XI0.XI1<9>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_61 XI1.XI0.XI1<9>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_66 XI1.XI0.XI1<9>.XI7<6>.NET_003
+ XI1.XI0.XI1<9>.XI7<6>.NET_000 XI1.XI0.XI1<9>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_72 XI1.XI0.XI1<9>.XI7<6>.NET_007
+ XI1.XI0.XI1<9>.XI7<6>.NET_001 XI1.XI0.XI1<9>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<6>.NET_005
+ XI1.XI0.XI1<9>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<6>.NET_003
+ XI1.XI0.XI1<9>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_41_11 REG_DATA_9<5> XI1.XI0.XI1<9>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<5>.MM_i_7 XI1.XI0.XI1<9>.XI7<5>.NET_001
+ XI1.XI0.XI1<9>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_13 XI1.XI0.XI1<9>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_18 XI1.XI0.XI1<9>.XI7<5>.NET_003
+ XI1.XI0.XI1<9>.XI7<5>.NET_001 XI1.XI0.XI1<9>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_24 XI1.XI0.XI1<9>.XI7<5>.NET_004
+ XI1.XI0.XI1<9>.XI7<5>.NET_000 XI1.XI0.XI1<9>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<5>.NET_005
+ XI1.XI0.XI1<9>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<5>.NET_003
+ XI1.XI0.XI1<9>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_89_4 REG_DATA_9<5> XI1.XI0.XI1<9>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<5>.MM_i_55 XI1.XI0.XI1<9>.XI7<5>.NET_001
+ XI1.XI0.XI1<9>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_61 XI1.XI0.XI1<9>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_66 XI1.XI0.XI1<9>.XI7<5>.NET_003
+ XI1.XI0.XI1<9>.XI7<5>.NET_000 XI1.XI0.XI1<9>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_72 XI1.XI0.XI1<9>.XI7<5>.NET_007
+ XI1.XI0.XI1<9>.XI7<5>.NET_001 XI1.XI0.XI1<9>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<5>.NET_005
+ XI1.XI0.XI1<9>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<5>.NET_003
+ XI1.XI0.XI1<9>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_41_11 REG_DATA_9<4> XI1.XI0.XI1<9>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<4>.MM_i_7 XI1.XI0.XI1<9>.XI7<4>.NET_001
+ XI1.XI0.XI1<9>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_13 XI1.XI0.XI1<9>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_18 XI1.XI0.XI1<9>.XI7<4>.NET_003
+ XI1.XI0.XI1<9>.XI7<4>.NET_001 XI1.XI0.XI1<9>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_24 XI1.XI0.XI1<9>.XI7<4>.NET_004
+ XI1.XI0.XI1<9>.XI7<4>.NET_000 XI1.XI0.XI1<9>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<4>.NET_005
+ XI1.XI0.XI1<9>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<4>.NET_003
+ XI1.XI0.XI1<9>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_89_4 REG_DATA_9<4> XI1.XI0.XI1<9>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<4>.MM_i_55 XI1.XI0.XI1<9>.XI7<4>.NET_001
+ XI1.XI0.XI1<9>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_61 XI1.XI0.XI1<9>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_66 XI1.XI0.XI1<9>.XI7<4>.NET_003
+ XI1.XI0.XI1<9>.XI7<4>.NET_000 XI1.XI0.XI1<9>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_72 XI1.XI0.XI1<9>.XI7<4>.NET_007
+ XI1.XI0.XI1<9>.XI7<4>.NET_001 XI1.XI0.XI1<9>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<4>.NET_005
+ XI1.XI0.XI1<9>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<4>.NET_003
+ XI1.XI0.XI1<9>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_41_11 REG_DATA_9<11> XI1.XI0.XI1<9>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<11>.MM_i_7 XI1.XI0.XI1<9>.XI7<11>.NET_001
+ XI1.XI0.XI1<9>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_13 XI1.XI0.XI1<9>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_18 XI1.XI0.XI1<9>.XI7<11>.NET_003
+ XI1.XI0.XI1<9>.XI7<11>.NET_001 XI1.XI0.XI1<9>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_24 XI1.XI0.XI1<9>.XI7<11>.NET_004
+ XI1.XI0.XI1<9>.XI7<11>.NET_000 XI1.XI0.XI1<9>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<11>.NET_005
+ XI1.XI0.XI1<9>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<11>.NET_003
+ XI1.XI0.XI1<9>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_89_4 REG_DATA_9<11> XI1.XI0.XI1<9>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<11>.MM_i_55 XI1.XI0.XI1<9>.XI7<11>.NET_001
+ XI1.XI0.XI1<9>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_61 XI1.XI0.XI1<9>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_66 XI1.XI0.XI1<9>.XI7<11>.NET_003
+ XI1.XI0.XI1<9>.XI7<11>.NET_000 XI1.XI0.XI1<9>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_72 XI1.XI0.XI1<9>.XI7<11>.NET_007
+ XI1.XI0.XI1<9>.XI7<11>.NET_001 XI1.XI0.XI1<9>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<11>.NET_005
+ XI1.XI0.XI1<9>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<11>.NET_003
+ XI1.XI0.XI1<9>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_41_11 REG_DATA_9<10> XI1.XI0.XI1<9>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<10>.MM_i_7 XI1.XI0.XI1<9>.XI7<10>.NET_001
+ XI1.XI0.XI1<9>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_13 XI1.XI0.XI1<9>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_18 XI1.XI0.XI1<9>.XI7<10>.NET_003
+ XI1.XI0.XI1<9>.XI7<10>.NET_001 XI1.XI0.XI1<9>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_24 XI1.XI0.XI1<9>.XI7<10>.NET_004
+ XI1.XI0.XI1<9>.XI7<10>.NET_000 XI1.XI0.XI1<9>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<10>.NET_005
+ XI1.XI0.XI1<9>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<10>.NET_003
+ XI1.XI0.XI1<9>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_89_4 REG_DATA_9<10> XI1.XI0.XI1<9>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<10>.MM_i_55 XI1.XI0.XI1<9>.XI7<10>.NET_001
+ XI1.XI0.XI1<9>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_61 XI1.XI0.XI1<9>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_66 XI1.XI0.XI1<9>.XI7<10>.NET_003
+ XI1.XI0.XI1<9>.XI7<10>.NET_000 XI1.XI0.XI1<9>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_72 XI1.XI0.XI1<9>.XI7<10>.NET_007
+ XI1.XI0.XI1<9>.XI7<10>.NET_001 XI1.XI0.XI1<9>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<10>.NET_005
+ XI1.XI0.XI1<9>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<10>.NET_003
+ XI1.XI0.XI1<9>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_41_11 REG_DATA_9<9> XI1.XI0.XI1<9>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<9>.MM_i_7 XI1.XI0.XI1<9>.XI7<9>.NET_001
+ XI1.XI0.XI1<9>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_13 XI1.XI0.XI1<9>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_18 XI1.XI0.XI1<9>.XI7<9>.NET_003
+ XI1.XI0.XI1<9>.XI7<9>.NET_001 XI1.XI0.XI1<9>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_24 XI1.XI0.XI1<9>.XI7<9>.NET_004
+ XI1.XI0.XI1<9>.XI7<9>.NET_000 XI1.XI0.XI1<9>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<9>.NET_005
+ XI1.XI0.XI1<9>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<9>.NET_003
+ XI1.XI0.XI1<9>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_89_4 REG_DATA_9<9> XI1.XI0.XI1<9>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<9>.MM_i_55 XI1.XI0.XI1<9>.XI7<9>.NET_001
+ XI1.XI0.XI1<9>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_61 XI1.XI0.XI1<9>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_66 XI1.XI0.XI1<9>.XI7<9>.NET_003
+ XI1.XI0.XI1<9>.XI7<9>.NET_000 XI1.XI0.XI1<9>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_72 XI1.XI0.XI1<9>.XI7<9>.NET_007
+ XI1.XI0.XI1<9>.XI7<9>.NET_001 XI1.XI0.XI1<9>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<9>.NET_005
+ XI1.XI0.XI1<9>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<9>.NET_003
+ XI1.XI0.XI1<9>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_41_11 REG_DATA_9<8> XI1.XI0.XI1<9>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<8>.MM_i_7 XI1.XI0.XI1<9>.XI7<8>.NET_001
+ XI1.XI0.XI1<9>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_13 XI1.XI0.XI1<9>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_18 XI1.XI0.XI1<9>.XI7<8>.NET_003
+ XI1.XI0.XI1<9>.XI7<8>.NET_001 XI1.XI0.XI1<9>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_24 XI1.XI0.XI1<9>.XI7<8>.NET_004
+ XI1.XI0.XI1<9>.XI7<8>.NET_000 XI1.XI0.XI1<9>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<8>.NET_005
+ XI1.XI0.XI1<9>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<8>.NET_003
+ XI1.XI0.XI1<9>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_89_4 REG_DATA_9<8> XI1.XI0.XI1<9>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<8>.MM_i_55 XI1.XI0.XI1<9>.XI7<8>.NET_001
+ XI1.XI0.XI1<9>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_61 XI1.XI0.XI1<9>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_66 XI1.XI0.XI1<9>.XI7<8>.NET_003
+ XI1.XI0.XI1<9>.XI7<8>.NET_000 XI1.XI0.XI1<9>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_72 XI1.XI0.XI1<9>.XI7<8>.NET_007
+ XI1.XI0.XI1<9>.XI7<8>.NET_001 XI1.XI0.XI1<9>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<8>.NET_005
+ XI1.XI0.XI1<9>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<8>.NET_003
+ XI1.XI0.XI1<9>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_41_11 REG_DATA_9<15> XI1.XI0.XI1<9>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<15>.MM_i_7 XI1.XI0.XI1<9>.XI7<15>.NET_001
+ XI1.XI0.XI1<9>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_13 XI1.XI0.XI1<9>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_18 XI1.XI0.XI1<9>.XI7<15>.NET_003
+ XI1.XI0.XI1<9>.XI7<15>.NET_001 XI1.XI0.XI1<9>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_24 XI1.XI0.XI1<9>.XI7<15>.NET_004
+ XI1.XI0.XI1<9>.XI7<15>.NET_000 XI1.XI0.XI1<9>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<15>.NET_005
+ XI1.XI0.XI1<9>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<15>.NET_003
+ XI1.XI0.XI1<9>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_89_4 REG_DATA_9<15> XI1.XI0.XI1<9>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<15>.MM_i_55 XI1.XI0.XI1<9>.XI7<15>.NET_001
+ XI1.XI0.XI1<9>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_61 XI1.XI0.XI1<9>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_66 XI1.XI0.XI1<9>.XI7<15>.NET_003
+ XI1.XI0.XI1<9>.XI7<15>.NET_000 XI1.XI0.XI1<9>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_72 XI1.XI0.XI1<9>.XI7<15>.NET_007
+ XI1.XI0.XI1<9>.XI7<15>.NET_001 XI1.XI0.XI1<9>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<15>.NET_005
+ XI1.XI0.XI1<9>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<15>.NET_003
+ XI1.XI0.XI1<9>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_41_11 REG_DATA_9<14> XI1.XI0.XI1<9>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<14>.MM_i_7 XI1.XI0.XI1<9>.XI7<14>.NET_001
+ XI1.XI0.XI1<9>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_13 XI1.XI0.XI1<9>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_18 XI1.XI0.XI1<9>.XI7<14>.NET_003
+ XI1.XI0.XI1<9>.XI7<14>.NET_001 XI1.XI0.XI1<9>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_24 XI1.XI0.XI1<9>.XI7<14>.NET_004
+ XI1.XI0.XI1<9>.XI7<14>.NET_000 XI1.XI0.XI1<9>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<14>.NET_005
+ XI1.XI0.XI1<9>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<14>.NET_003
+ XI1.XI0.XI1<9>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_89_4 REG_DATA_9<14> XI1.XI0.XI1<9>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<14>.MM_i_55 XI1.XI0.XI1<9>.XI7<14>.NET_001
+ XI1.XI0.XI1<9>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_61 XI1.XI0.XI1<9>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_66 XI1.XI0.XI1<9>.XI7<14>.NET_003
+ XI1.XI0.XI1<9>.XI7<14>.NET_000 XI1.XI0.XI1<9>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_72 XI1.XI0.XI1<9>.XI7<14>.NET_007
+ XI1.XI0.XI1<9>.XI7<14>.NET_001 XI1.XI0.XI1<9>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<14>.NET_005
+ XI1.XI0.XI1<9>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<14>.NET_003
+ XI1.XI0.XI1<9>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_41_11 REG_DATA_9<13> XI1.XI0.XI1<9>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<13>.MM_i_7 XI1.XI0.XI1<9>.XI7<13>.NET_001
+ XI1.XI0.XI1<9>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_13 XI1.XI0.XI1<9>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_18 XI1.XI0.XI1<9>.XI7<13>.NET_003
+ XI1.XI0.XI1<9>.XI7<13>.NET_001 XI1.XI0.XI1<9>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_24 XI1.XI0.XI1<9>.XI7<13>.NET_004
+ XI1.XI0.XI1<9>.XI7<13>.NET_000 XI1.XI0.XI1<9>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<13>.NET_005
+ XI1.XI0.XI1<9>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<13>.NET_003
+ XI1.XI0.XI1<9>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_89_4 REG_DATA_9<13> XI1.XI0.XI1<9>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<13>.MM_i_55 XI1.XI0.XI1<9>.XI7<13>.NET_001
+ XI1.XI0.XI1<9>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_61 XI1.XI0.XI1<9>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_66 XI1.XI0.XI1<9>.XI7<13>.NET_003
+ XI1.XI0.XI1<9>.XI7<13>.NET_000 XI1.XI0.XI1<9>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_72 XI1.XI0.XI1<9>.XI7<13>.NET_007
+ XI1.XI0.XI1<9>.XI7<13>.NET_001 XI1.XI0.XI1<9>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<13>.NET_005
+ XI1.XI0.XI1<9>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<13>.NET_003
+ XI1.XI0.XI1<9>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_41_11 REG_DATA_9<12> XI1.XI0.XI1<9>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<9>.XI7<12>.MM_i_7 XI1.XI0.XI1<9>.XI7<12>.NET_001
+ XI1.XI0.XI1<9>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_13 XI1.XI0.XI1<9>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_18 XI1.XI0.XI1<9>.XI7<12>.NET_003
+ XI1.XI0.XI1<9>.XI7<12>.NET_001 XI1.XI0.XI1<9>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_24 XI1.XI0.XI1<9>.XI7<12>.NET_004
+ XI1.XI0.XI1<9>.XI7<12>.NET_000 XI1.XI0.XI1<9>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<9>.XI7<12>.NET_005
+ XI1.XI0.XI1<9>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<9>.XI7<12>.NET_003
+ XI1.XI0.XI1<9>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<9>
+ XI1.XI0.XI1<9>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_89_4 REG_DATA_9<12> XI1.XI0.XI1<9>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<9>.XI7<12>.MM_i_55 XI1.XI0.XI1<9>.XI7<12>.NET_001
+ XI1.XI0.XI1<9>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_61 XI1.XI0.XI1<9>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_66 XI1.XI0.XI1<9>.XI7<12>.NET_003
+ XI1.XI0.XI1<9>.XI7<12>.NET_000 XI1.XI0.XI1<9>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_72 XI1.XI0.XI1<9>.XI7<12>.NET_007
+ XI1.XI0.XI1<9>.XI7<12>.NET_001 XI1.XI0.XI1<9>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<9>.XI7<12>.NET_005
+ XI1.XI0.XI1<9>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<9>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<9>.XI7<12>.NET_003
+ XI1.XI0.XI1<9>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_41_11 REG_DATA_8<3> XI1.XI0.XI1<8>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<3>.MM_i_7 XI1.XI0.XI1<8>.XI7<3>.NET_001
+ XI1.XI0.XI1<8>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_13 XI1.XI0.XI1<8>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_18 XI1.XI0.XI1<8>.XI7<3>.NET_003
+ XI1.XI0.XI1<8>.XI7<3>.NET_001 XI1.XI0.XI1<8>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_24 XI1.XI0.XI1<8>.XI7<3>.NET_004
+ XI1.XI0.XI1<8>.XI7<3>.NET_000 XI1.XI0.XI1<8>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<3>.NET_005
+ XI1.XI0.XI1<8>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<3>.NET_003
+ XI1.XI0.XI1<8>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_89_4 REG_DATA_8<3> XI1.XI0.XI1<8>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<3>.MM_i_55 XI1.XI0.XI1<8>.XI7<3>.NET_001
+ XI1.XI0.XI1<8>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_61 XI1.XI0.XI1<8>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_66 XI1.XI0.XI1<8>.XI7<3>.NET_003
+ XI1.XI0.XI1<8>.XI7<3>.NET_000 XI1.XI0.XI1<8>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_72 XI1.XI0.XI1<8>.XI7<3>.NET_007
+ XI1.XI0.XI1<8>.XI7<3>.NET_001 XI1.XI0.XI1<8>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<3>.NET_005
+ XI1.XI0.XI1<8>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<3>.NET_003
+ XI1.XI0.XI1<8>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_41_11 REG_DATA_8<2> XI1.XI0.XI1<8>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<2>.MM_i_7 XI1.XI0.XI1<8>.XI7<2>.NET_001
+ XI1.XI0.XI1<8>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_13 XI1.XI0.XI1<8>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_18 XI1.XI0.XI1<8>.XI7<2>.NET_003
+ XI1.XI0.XI1<8>.XI7<2>.NET_001 XI1.XI0.XI1<8>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_24 XI1.XI0.XI1<8>.XI7<2>.NET_004
+ XI1.XI0.XI1<8>.XI7<2>.NET_000 XI1.XI0.XI1<8>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<2>.NET_005
+ XI1.XI0.XI1<8>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<2>.NET_003
+ XI1.XI0.XI1<8>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_89_4 REG_DATA_8<2> XI1.XI0.XI1<8>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<2>.MM_i_55 XI1.XI0.XI1<8>.XI7<2>.NET_001
+ XI1.XI0.XI1<8>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_61 XI1.XI0.XI1<8>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_66 XI1.XI0.XI1<8>.XI7<2>.NET_003
+ XI1.XI0.XI1<8>.XI7<2>.NET_000 XI1.XI0.XI1<8>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_72 XI1.XI0.XI1<8>.XI7<2>.NET_007
+ XI1.XI0.XI1<8>.XI7<2>.NET_001 XI1.XI0.XI1<8>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<2>.NET_005
+ XI1.XI0.XI1<8>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<2>.NET_003
+ XI1.XI0.XI1<8>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_41_11 REG_DATA_8<1> XI1.XI0.XI1<8>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<1>.MM_i_7 XI1.XI0.XI1<8>.XI7<1>.NET_001
+ XI1.XI0.XI1<8>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_13 XI1.XI0.XI1<8>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_18 XI1.XI0.XI1<8>.XI7<1>.NET_003
+ XI1.XI0.XI1<8>.XI7<1>.NET_001 XI1.XI0.XI1<8>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_24 XI1.XI0.XI1<8>.XI7<1>.NET_004
+ XI1.XI0.XI1<8>.XI7<1>.NET_000 XI1.XI0.XI1<8>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<1>.NET_005
+ XI1.XI0.XI1<8>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<1>.NET_003
+ XI1.XI0.XI1<8>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_89_4 REG_DATA_8<1> XI1.XI0.XI1<8>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<1>.MM_i_55 XI1.XI0.XI1<8>.XI7<1>.NET_001
+ XI1.XI0.XI1<8>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_61 XI1.XI0.XI1<8>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_66 XI1.XI0.XI1<8>.XI7<1>.NET_003
+ XI1.XI0.XI1<8>.XI7<1>.NET_000 XI1.XI0.XI1<8>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_72 XI1.XI0.XI1<8>.XI7<1>.NET_007
+ XI1.XI0.XI1<8>.XI7<1>.NET_001 XI1.XI0.XI1<8>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<1>.NET_005
+ XI1.XI0.XI1<8>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<1>.NET_003
+ XI1.XI0.XI1<8>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_41_11 REG_DATA_8<0> XI1.XI0.XI1<8>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<0>.MM_i_7 XI1.XI0.XI1<8>.XI7<0>.NET_001
+ XI1.XI0.XI1<8>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_13 XI1.XI0.XI1<8>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_18 XI1.XI0.XI1<8>.XI7<0>.NET_003
+ XI1.XI0.XI1<8>.XI7<0>.NET_001 XI1.XI0.XI1<8>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_24 XI1.XI0.XI1<8>.XI7<0>.NET_004
+ XI1.XI0.XI1<8>.XI7<0>.NET_000 XI1.XI0.XI1<8>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<0>.NET_005
+ XI1.XI0.XI1<8>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<0>.NET_003
+ XI1.XI0.XI1<8>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_89_4 REG_DATA_8<0> XI1.XI0.XI1<8>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<0>.MM_i_55 XI1.XI0.XI1<8>.XI7<0>.NET_001
+ XI1.XI0.XI1<8>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_61 XI1.XI0.XI1<8>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_66 XI1.XI0.XI1<8>.XI7<0>.NET_003
+ XI1.XI0.XI1<8>.XI7<0>.NET_000 XI1.XI0.XI1<8>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_72 XI1.XI0.XI1<8>.XI7<0>.NET_007
+ XI1.XI0.XI1<8>.XI7<0>.NET_001 XI1.XI0.XI1<8>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<0>.NET_005
+ XI1.XI0.XI1<8>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<0>.NET_003
+ XI1.XI0.XI1<8>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_41_11 REG_DATA_8<7> XI1.XI0.XI1<8>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<7>.MM_i_7 XI1.XI0.XI1<8>.XI7<7>.NET_001
+ XI1.XI0.XI1<8>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_13 XI1.XI0.XI1<8>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_18 XI1.XI0.XI1<8>.XI7<7>.NET_003
+ XI1.XI0.XI1<8>.XI7<7>.NET_001 XI1.XI0.XI1<8>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_24 XI1.XI0.XI1<8>.XI7<7>.NET_004
+ XI1.XI0.XI1<8>.XI7<7>.NET_000 XI1.XI0.XI1<8>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<7>.NET_005
+ XI1.XI0.XI1<8>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<7>.NET_003
+ XI1.XI0.XI1<8>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_89_4 REG_DATA_8<7> XI1.XI0.XI1<8>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<7>.MM_i_55 XI1.XI0.XI1<8>.XI7<7>.NET_001
+ XI1.XI0.XI1<8>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_61 XI1.XI0.XI1<8>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_66 XI1.XI0.XI1<8>.XI7<7>.NET_003
+ XI1.XI0.XI1<8>.XI7<7>.NET_000 XI1.XI0.XI1<8>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_72 XI1.XI0.XI1<8>.XI7<7>.NET_007
+ XI1.XI0.XI1<8>.XI7<7>.NET_001 XI1.XI0.XI1<8>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<7>.NET_005
+ XI1.XI0.XI1<8>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<7>.NET_003
+ XI1.XI0.XI1<8>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_41_11 REG_DATA_8<6> XI1.XI0.XI1<8>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<6>.MM_i_7 XI1.XI0.XI1<8>.XI7<6>.NET_001
+ XI1.XI0.XI1<8>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_13 XI1.XI0.XI1<8>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_18 XI1.XI0.XI1<8>.XI7<6>.NET_003
+ XI1.XI0.XI1<8>.XI7<6>.NET_001 XI1.XI0.XI1<8>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_24 XI1.XI0.XI1<8>.XI7<6>.NET_004
+ XI1.XI0.XI1<8>.XI7<6>.NET_000 XI1.XI0.XI1<8>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<6>.NET_005
+ XI1.XI0.XI1<8>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<6>.NET_003
+ XI1.XI0.XI1<8>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_89_4 REG_DATA_8<6> XI1.XI0.XI1<8>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<6>.MM_i_55 XI1.XI0.XI1<8>.XI7<6>.NET_001
+ XI1.XI0.XI1<8>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_61 XI1.XI0.XI1<8>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_66 XI1.XI0.XI1<8>.XI7<6>.NET_003
+ XI1.XI0.XI1<8>.XI7<6>.NET_000 XI1.XI0.XI1<8>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_72 XI1.XI0.XI1<8>.XI7<6>.NET_007
+ XI1.XI0.XI1<8>.XI7<6>.NET_001 XI1.XI0.XI1<8>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<6>.NET_005
+ XI1.XI0.XI1<8>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<6>.NET_003
+ XI1.XI0.XI1<8>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_41_11 REG_DATA_8<5> XI1.XI0.XI1<8>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<5>.MM_i_7 XI1.XI0.XI1<8>.XI7<5>.NET_001
+ XI1.XI0.XI1<8>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_13 XI1.XI0.XI1<8>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_18 XI1.XI0.XI1<8>.XI7<5>.NET_003
+ XI1.XI0.XI1<8>.XI7<5>.NET_001 XI1.XI0.XI1<8>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_24 XI1.XI0.XI1<8>.XI7<5>.NET_004
+ XI1.XI0.XI1<8>.XI7<5>.NET_000 XI1.XI0.XI1<8>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<5>.NET_005
+ XI1.XI0.XI1<8>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<5>.NET_003
+ XI1.XI0.XI1<8>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_89_4 REG_DATA_8<5> XI1.XI0.XI1<8>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<5>.MM_i_55 XI1.XI0.XI1<8>.XI7<5>.NET_001
+ XI1.XI0.XI1<8>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_61 XI1.XI0.XI1<8>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_66 XI1.XI0.XI1<8>.XI7<5>.NET_003
+ XI1.XI0.XI1<8>.XI7<5>.NET_000 XI1.XI0.XI1<8>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_72 XI1.XI0.XI1<8>.XI7<5>.NET_007
+ XI1.XI0.XI1<8>.XI7<5>.NET_001 XI1.XI0.XI1<8>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<5>.NET_005
+ XI1.XI0.XI1<8>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<5>.NET_003
+ XI1.XI0.XI1<8>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_41_11 REG_DATA_8<4> XI1.XI0.XI1<8>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<4>.MM_i_7 XI1.XI0.XI1<8>.XI7<4>.NET_001
+ XI1.XI0.XI1<8>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_13 XI1.XI0.XI1<8>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_18 XI1.XI0.XI1<8>.XI7<4>.NET_003
+ XI1.XI0.XI1<8>.XI7<4>.NET_001 XI1.XI0.XI1<8>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_24 XI1.XI0.XI1<8>.XI7<4>.NET_004
+ XI1.XI0.XI1<8>.XI7<4>.NET_000 XI1.XI0.XI1<8>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<4>.NET_005
+ XI1.XI0.XI1<8>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<4>.NET_003
+ XI1.XI0.XI1<8>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_89_4 REG_DATA_8<4> XI1.XI0.XI1<8>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<4>.MM_i_55 XI1.XI0.XI1<8>.XI7<4>.NET_001
+ XI1.XI0.XI1<8>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_61 XI1.XI0.XI1<8>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_66 XI1.XI0.XI1<8>.XI7<4>.NET_003
+ XI1.XI0.XI1<8>.XI7<4>.NET_000 XI1.XI0.XI1<8>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_72 XI1.XI0.XI1<8>.XI7<4>.NET_007
+ XI1.XI0.XI1<8>.XI7<4>.NET_001 XI1.XI0.XI1<8>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<4>.NET_005
+ XI1.XI0.XI1<8>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<4>.NET_003
+ XI1.XI0.XI1<8>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_41_11 REG_DATA_8<11> XI1.XI0.XI1<8>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<11>.MM_i_7 XI1.XI0.XI1<8>.XI7<11>.NET_001
+ XI1.XI0.XI1<8>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_13 XI1.XI0.XI1<8>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_18 XI1.XI0.XI1<8>.XI7<11>.NET_003
+ XI1.XI0.XI1<8>.XI7<11>.NET_001 XI1.XI0.XI1<8>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_24 XI1.XI0.XI1<8>.XI7<11>.NET_004
+ XI1.XI0.XI1<8>.XI7<11>.NET_000 XI1.XI0.XI1<8>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<11>.NET_005
+ XI1.XI0.XI1<8>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<11>.NET_003
+ XI1.XI0.XI1<8>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_89_4 REG_DATA_8<11> XI1.XI0.XI1<8>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<11>.MM_i_55 XI1.XI0.XI1<8>.XI7<11>.NET_001
+ XI1.XI0.XI1<8>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_61 XI1.XI0.XI1<8>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_66 XI1.XI0.XI1<8>.XI7<11>.NET_003
+ XI1.XI0.XI1<8>.XI7<11>.NET_000 XI1.XI0.XI1<8>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_72 XI1.XI0.XI1<8>.XI7<11>.NET_007
+ XI1.XI0.XI1<8>.XI7<11>.NET_001 XI1.XI0.XI1<8>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<11>.NET_005
+ XI1.XI0.XI1<8>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<11>.NET_003
+ XI1.XI0.XI1<8>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_41_11 REG_DATA_8<10> XI1.XI0.XI1<8>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<10>.MM_i_7 XI1.XI0.XI1<8>.XI7<10>.NET_001
+ XI1.XI0.XI1<8>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_13 XI1.XI0.XI1<8>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_18 XI1.XI0.XI1<8>.XI7<10>.NET_003
+ XI1.XI0.XI1<8>.XI7<10>.NET_001 XI1.XI0.XI1<8>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_24 XI1.XI0.XI1<8>.XI7<10>.NET_004
+ XI1.XI0.XI1<8>.XI7<10>.NET_000 XI1.XI0.XI1<8>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<10>.NET_005
+ XI1.XI0.XI1<8>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<10>.NET_003
+ XI1.XI0.XI1<8>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_89_4 REG_DATA_8<10> XI1.XI0.XI1<8>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<10>.MM_i_55 XI1.XI0.XI1<8>.XI7<10>.NET_001
+ XI1.XI0.XI1<8>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_61 XI1.XI0.XI1<8>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_66 XI1.XI0.XI1<8>.XI7<10>.NET_003
+ XI1.XI0.XI1<8>.XI7<10>.NET_000 XI1.XI0.XI1<8>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_72 XI1.XI0.XI1<8>.XI7<10>.NET_007
+ XI1.XI0.XI1<8>.XI7<10>.NET_001 XI1.XI0.XI1<8>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<10>.NET_005
+ XI1.XI0.XI1<8>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<10>.NET_003
+ XI1.XI0.XI1<8>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_41_11 REG_DATA_8<9> XI1.XI0.XI1<8>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<9>.MM_i_7 XI1.XI0.XI1<8>.XI7<9>.NET_001
+ XI1.XI0.XI1<8>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_13 XI1.XI0.XI1<8>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_18 XI1.XI0.XI1<8>.XI7<9>.NET_003
+ XI1.XI0.XI1<8>.XI7<9>.NET_001 XI1.XI0.XI1<8>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_24 XI1.XI0.XI1<8>.XI7<9>.NET_004
+ XI1.XI0.XI1<8>.XI7<9>.NET_000 XI1.XI0.XI1<8>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<9>.NET_005
+ XI1.XI0.XI1<8>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<9>.NET_003
+ XI1.XI0.XI1<8>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_89_4 REG_DATA_8<9> XI1.XI0.XI1<8>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<9>.MM_i_55 XI1.XI0.XI1<8>.XI7<9>.NET_001
+ XI1.XI0.XI1<8>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_61 XI1.XI0.XI1<8>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_66 XI1.XI0.XI1<8>.XI7<9>.NET_003
+ XI1.XI0.XI1<8>.XI7<9>.NET_000 XI1.XI0.XI1<8>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_72 XI1.XI0.XI1<8>.XI7<9>.NET_007
+ XI1.XI0.XI1<8>.XI7<9>.NET_001 XI1.XI0.XI1<8>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<9>.NET_005
+ XI1.XI0.XI1<8>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<9>.NET_003
+ XI1.XI0.XI1<8>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_41_11 REG_DATA_8<8> XI1.XI0.XI1<8>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<8>.MM_i_7 XI1.XI0.XI1<8>.XI7<8>.NET_001
+ XI1.XI0.XI1<8>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_13 XI1.XI0.XI1<8>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_18 XI1.XI0.XI1<8>.XI7<8>.NET_003
+ XI1.XI0.XI1<8>.XI7<8>.NET_001 XI1.XI0.XI1<8>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_24 XI1.XI0.XI1<8>.XI7<8>.NET_004
+ XI1.XI0.XI1<8>.XI7<8>.NET_000 XI1.XI0.XI1<8>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<8>.NET_005
+ XI1.XI0.XI1<8>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<8>.NET_003
+ XI1.XI0.XI1<8>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_89_4 REG_DATA_8<8> XI1.XI0.XI1<8>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<8>.MM_i_55 XI1.XI0.XI1<8>.XI7<8>.NET_001
+ XI1.XI0.XI1<8>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_61 XI1.XI0.XI1<8>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_66 XI1.XI0.XI1<8>.XI7<8>.NET_003
+ XI1.XI0.XI1<8>.XI7<8>.NET_000 XI1.XI0.XI1<8>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_72 XI1.XI0.XI1<8>.XI7<8>.NET_007
+ XI1.XI0.XI1<8>.XI7<8>.NET_001 XI1.XI0.XI1<8>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<8>.NET_005
+ XI1.XI0.XI1<8>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<8>.NET_003
+ XI1.XI0.XI1<8>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_41_11 REG_DATA_8<15> XI1.XI0.XI1<8>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<15>.MM_i_7 XI1.XI0.XI1<8>.XI7<15>.NET_001
+ XI1.XI0.XI1<8>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_13 XI1.XI0.XI1<8>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_18 XI1.XI0.XI1<8>.XI7<15>.NET_003
+ XI1.XI0.XI1<8>.XI7<15>.NET_001 XI1.XI0.XI1<8>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_24 XI1.XI0.XI1<8>.XI7<15>.NET_004
+ XI1.XI0.XI1<8>.XI7<15>.NET_000 XI1.XI0.XI1<8>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<15>.NET_005
+ XI1.XI0.XI1<8>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<15>.NET_003
+ XI1.XI0.XI1<8>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_89_4 REG_DATA_8<15> XI1.XI0.XI1<8>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<15>.MM_i_55 XI1.XI0.XI1<8>.XI7<15>.NET_001
+ XI1.XI0.XI1<8>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_61 XI1.XI0.XI1<8>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_66 XI1.XI0.XI1<8>.XI7<15>.NET_003
+ XI1.XI0.XI1<8>.XI7<15>.NET_000 XI1.XI0.XI1<8>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_72 XI1.XI0.XI1<8>.XI7<15>.NET_007
+ XI1.XI0.XI1<8>.XI7<15>.NET_001 XI1.XI0.XI1<8>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<15>.NET_005
+ XI1.XI0.XI1<8>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<15>.NET_003
+ XI1.XI0.XI1<8>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_41_11 REG_DATA_8<14> XI1.XI0.XI1<8>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<14>.MM_i_7 XI1.XI0.XI1<8>.XI7<14>.NET_001
+ XI1.XI0.XI1<8>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_13 XI1.XI0.XI1<8>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_18 XI1.XI0.XI1<8>.XI7<14>.NET_003
+ XI1.XI0.XI1<8>.XI7<14>.NET_001 XI1.XI0.XI1<8>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_24 XI1.XI0.XI1<8>.XI7<14>.NET_004
+ XI1.XI0.XI1<8>.XI7<14>.NET_000 XI1.XI0.XI1<8>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<14>.NET_005
+ XI1.XI0.XI1<8>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<14>.NET_003
+ XI1.XI0.XI1<8>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_89_4 REG_DATA_8<14> XI1.XI0.XI1<8>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<14>.MM_i_55 XI1.XI0.XI1<8>.XI7<14>.NET_001
+ XI1.XI0.XI1<8>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_61 XI1.XI0.XI1<8>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_66 XI1.XI0.XI1<8>.XI7<14>.NET_003
+ XI1.XI0.XI1<8>.XI7<14>.NET_000 XI1.XI0.XI1<8>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_72 XI1.XI0.XI1<8>.XI7<14>.NET_007
+ XI1.XI0.XI1<8>.XI7<14>.NET_001 XI1.XI0.XI1<8>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<14>.NET_005
+ XI1.XI0.XI1<8>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<14>.NET_003
+ XI1.XI0.XI1<8>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_41_11 REG_DATA_8<13> XI1.XI0.XI1<8>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<13>.MM_i_7 XI1.XI0.XI1<8>.XI7<13>.NET_001
+ XI1.XI0.XI1<8>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_13 XI1.XI0.XI1<8>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_18 XI1.XI0.XI1<8>.XI7<13>.NET_003
+ XI1.XI0.XI1<8>.XI7<13>.NET_001 XI1.XI0.XI1<8>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_24 XI1.XI0.XI1<8>.XI7<13>.NET_004
+ XI1.XI0.XI1<8>.XI7<13>.NET_000 XI1.XI0.XI1<8>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<13>.NET_005
+ XI1.XI0.XI1<8>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<13>.NET_003
+ XI1.XI0.XI1<8>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_89_4 REG_DATA_8<13> XI1.XI0.XI1<8>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<13>.MM_i_55 XI1.XI0.XI1<8>.XI7<13>.NET_001
+ XI1.XI0.XI1<8>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_61 XI1.XI0.XI1<8>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_66 XI1.XI0.XI1<8>.XI7<13>.NET_003
+ XI1.XI0.XI1<8>.XI7<13>.NET_000 XI1.XI0.XI1<8>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_72 XI1.XI0.XI1<8>.XI7<13>.NET_007
+ XI1.XI0.XI1<8>.XI7<13>.NET_001 XI1.XI0.XI1<8>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<13>.NET_005
+ XI1.XI0.XI1<8>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<13>.NET_003
+ XI1.XI0.XI1<8>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_41_11 REG_DATA_8<12> XI1.XI0.XI1<8>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<8>.XI7<12>.MM_i_7 XI1.XI0.XI1<8>.XI7<12>.NET_001
+ XI1.XI0.XI1<8>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_13 XI1.XI0.XI1<8>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_18 XI1.XI0.XI1<8>.XI7<12>.NET_003
+ XI1.XI0.XI1<8>.XI7<12>.NET_001 XI1.XI0.XI1<8>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_24 XI1.XI0.XI1<8>.XI7<12>.NET_004
+ XI1.XI0.XI1<8>.XI7<12>.NET_000 XI1.XI0.XI1<8>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<8>.XI7<12>.NET_005
+ XI1.XI0.XI1<8>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<8>.XI7<12>.NET_003
+ XI1.XI0.XI1<8>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<8>
+ XI1.XI0.XI1<8>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_89_4 REG_DATA_8<12> XI1.XI0.XI1<8>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<8>.XI7<12>.MM_i_55 XI1.XI0.XI1<8>.XI7<12>.NET_001
+ XI1.XI0.XI1<8>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_61 XI1.XI0.XI1<8>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_66 XI1.XI0.XI1<8>.XI7<12>.NET_003
+ XI1.XI0.XI1<8>.XI7<12>.NET_000 XI1.XI0.XI1<8>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_72 XI1.XI0.XI1<8>.XI7<12>.NET_007
+ XI1.XI0.XI1<8>.XI7<12>.NET_001 XI1.XI0.XI1<8>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<8>.XI7<12>.NET_005
+ XI1.XI0.XI1<8>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<8>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<8>.XI7<12>.NET_003
+ XI1.XI0.XI1<8>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_41_11 REG_DATA_7<3> XI1.XI0.XI1<7>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<3>.MM_i_7 XI1.XI0.XI1<7>.XI7<3>.NET_001
+ XI1.XI0.XI1<7>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_13 XI1.XI0.XI1<7>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_18 XI1.XI0.XI1<7>.XI7<3>.NET_003
+ XI1.XI0.XI1<7>.XI7<3>.NET_001 XI1.XI0.XI1<7>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_24 XI1.XI0.XI1<7>.XI7<3>.NET_004
+ XI1.XI0.XI1<7>.XI7<3>.NET_000 XI1.XI0.XI1<7>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<3>.NET_005
+ XI1.XI0.XI1<7>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<3>.NET_003
+ XI1.XI0.XI1<7>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_89_4 REG_DATA_7<3> XI1.XI0.XI1<7>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<3>.MM_i_55 XI1.XI0.XI1<7>.XI7<3>.NET_001
+ XI1.XI0.XI1<7>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_61 XI1.XI0.XI1<7>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_66 XI1.XI0.XI1<7>.XI7<3>.NET_003
+ XI1.XI0.XI1<7>.XI7<3>.NET_000 XI1.XI0.XI1<7>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_72 XI1.XI0.XI1<7>.XI7<3>.NET_007
+ XI1.XI0.XI1<7>.XI7<3>.NET_001 XI1.XI0.XI1<7>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<3>.NET_005
+ XI1.XI0.XI1<7>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<3>.NET_003
+ XI1.XI0.XI1<7>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_41_11 REG_DATA_7<2> XI1.XI0.XI1<7>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<2>.MM_i_7 XI1.XI0.XI1<7>.XI7<2>.NET_001
+ XI1.XI0.XI1<7>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_13 XI1.XI0.XI1<7>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_18 XI1.XI0.XI1<7>.XI7<2>.NET_003
+ XI1.XI0.XI1<7>.XI7<2>.NET_001 XI1.XI0.XI1<7>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_24 XI1.XI0.XI1<7>.XI7<2>.NET_004
+ XI1.XI0.XI1<7>.XI7<2>.NET_000 XI1.XI0.XI1<7>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<2>.NET_005
+ XI1.XI0.XI1<7>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<2>.NET_003
+ XI1.XI0.XI1<7>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_89_4 REG_DATA_7<2> XI1.XI0.XI1<7>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<2>.MM_i_55 XI1.XI0.XI1<7>.XI7<2>.NET_001
+ XI1.XI0.XI1<7>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_61 XI1.XI0.XI1<7>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_66 XI1.XI0.XI1<7>.XI7<2>.NET_003
+ XI1.XI0.XI1<7>.XI7<2>.NET_000 XI1.XI0.XI1<7>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_72 XI1.XI0.XI1<7>.XI7<2>.NET_007
+ XI1.XI0.XI1<7>.XI7<2>.NET_001 XI1.XI0.XI1<7>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<2>.NET_005
+ XI1.XI0.XI1<7>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<2>.NET_003
+ XI1.XI0.XI1<7>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_41_11 REG_DATA_7<1> XI1.XI0.XI1<7>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<1>.MM_i_7 XI1.XI0.XI1<7>.XI7<1>.NET_001
+ XI1.XI0.XI1<7>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_13 XI1.XI0.XI1<7>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_18 XI1.XI0.XI1<7>.XI7<1>.NET_003
+ XI1.XI0.XI1<7>.XI7<1>.NET_001 XI1.XI0.XI1<7>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_24 XI1.XI0.XI1<7>.XI7<1>.NET_004
+ XI1.XI0.XI1<7>.XI7<1>.NET_000 XI1.XI0.XI1<7>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<1>.NET_005
+ XI1.XI0.XI1<7>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<1>.NET_003
+ XI1.XI0.XI1<7>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_89_4 REG_DATA_7<1> XI1.XI0.XI1<7>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<1>.MM_i_55 XI1.XI0.XI1<7>.XI7<1>.NET_001
+ XI1.XI0.XI1<7>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_61 XI1.XI0.XI1<7>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_66 XI1.XI0.XI1<7>.XI7<1>.NET_003
+ XI1.XI0.XI1<7>.XI7<1>.NET_000 XI1.XI0.XI1<7>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_72 XI1.XI0.XI1<7>.XI7<1>.NET_007
+ XI1.XI0.XI1<7>.XI7<1>.NET_001 XI1.XI0.XI1<7>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<1>.NET_005
+ XI1.XI0.XI1<7>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<1>.NET_003
+ XI1.XI0.XI1<7>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_41_11 REG_DATA_7<0> XI1.XI0.XI1<7>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<0>.MM_i_7 XI1.XI0.XI1<7>.XI7<0>.NET_001
+ XI1.XI0.XI1<7>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_13 XI1.XI0.XI1<7>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_18 XI1.XI0.XI1<7>.XI7<0>.NET_003
+ XI1.XI0.XI1<7>.XI7<0>.NET_001 XI1.XI0.XI1<7>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_24 XI1.XI0.XI1<7>.XI7<0>.NET_004
+ XI1.XI0.XI1<7>.XI7<0>.NET_000 XI1.XI0.XI1<7>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<0>.NET_005
+ XI1.XI0.XI1<7>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<0>.NET_003
+ XI1.XI0.XI1<7>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_89_4 REG_DATA_7<0> XI1.XI0.XI1<7>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<0>.MM_i_55 XI1.XI0.XI1<7>.XI7<0>.NET_001
+ XI1.XI0.XI1<7>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_61 XI1.XI0.XI1<7>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_66 XI1.XI0.XI1<7>.XI7<0>.NET_003
+ XI1.XI0.XI1<7>.XI7<0>.NET_000 XI1.XI0.XI1<7>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_72 XI1.XI0.XI1<7>.XI7<0>.NET_007
+ XI1.XI0.XI1<7>.XI7<0>.NET_001 XI1.XI0.XI1<7>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<0>.NET_005
+ XI1.XI0.XI1<7>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<0>.NET_003
+ XI1.XI0.XI1<7>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_41_11 REG_DATA_7<7> XI1.XI0.XI1<7>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<7>.MM_i_7 XI1.XI0.XI1<7>.XI7<7>.NET_001
+ XI1.XI0.XI1<7>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_13 XI1.XI0.XI1<7>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_18 XI1.XI0.XI1<7>.XI7<7>.NET_003
+ XI1.XI0.XI1<7>.XI7<7>.NET_001 XI1.XI0.XI1<7>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_24 XI1.XI0.XI1<7>.XI7<7>.NET_004
+ XI1.XI0.XI1<7>.XI7<7>.NET_000 XI1.XI0.XI1<7>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<7>.NET_005
+ XI1.XI0.XI1<7>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<7>.NET_003
+ XI1.XI0.XI1<7>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_89_4 REG_DATA_7<7> XI1.XI0.XI1<7>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<7>.MM_i_55 XI1.XI0.XI1<7>.XI7<7>.NET_001
+ XI1.XI0.XI1<7>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_61 XI1.XI0.XI1<7>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_66 XI1.XI0.XI1<7>.XI7<7>.NET_003
+ XI1.XI0.XI1<7>.XI7<7>.NET_000 XI1.XI0.XI1<7>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_72 XI1.XI0.XI1<7>.XI7<7>.NET_007
+ XI1.XI0.XI1<7>.XI7<7>.NET_001 XI1.XI0.XI1<7>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<7>.NET_005
+ XI1.XI0.XI1<7>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<7>.NET_003
+ XI1.XI0.XI1<7>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_41_11 REG_DATA_7<6> XI1.XI0.XI1<7>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<6>.MM_i_7 XI1.XI0.XI1<7>.XI7<6>.NET_001
+ XI1.XI0.XI1<7>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_13 XI1.XI0.XI1<7>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_18 XI1.XI0.XI1<7>.XI7<6>.NET_003
+ XI1.XI0.XI1<7>.XI7<6>.NET_001 XI1.XI0.XI1<7>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_24 XI1.XI0.XI1<7>.XI7<6>.NET_004
+ XI1.XI0.XI1<7>.XI7<6>.NET_000 XI1.XI0.XI1<7>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<6>.NET_005
+ XI1.XI0.XI1<7>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<6>.NET_003
+ XI1.XI0.XI1<7>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_89_4 REG_DATA_7<6> XI1.XI0.XI1<7>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<6>.MM_i_55 XI1.XI0.XI1<7>.XI7<6>.NET_001
+ XI1.XI0.XI1<7>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_61 XI1.XI0.XI1<7>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_66 XI1.XI0.XI1<7>.XI7<6>.NET_003
+ XI1.XI0.XI1<7>.XI7<6>.NET_000 XI1.XI0.XI1<7>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_72 XI1.XI0.XI1<7>.XI7<6>.NET_007
+ XI1.XI0.XI1<7>.XI7<6>.NET_001 XI1.XI0.XI1<7>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<6>.NET_005
+ XI1.XI0.XI1<7>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<6>.NET_003
+ XI1.XI0.XI1<7>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_41_11 REG_DATA_7<5> XI1.XI0.XI1<7>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<5>.MM_i_7 XI1.XI0.XI1<7>.XI7<5>.NET_001
+ XI1.XI0.XI1<7>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_13 XI1.XI0.XI1<7>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_18 XI1.XI0.XI1<7>.XI7<5>.NET_003
+ XI1.XI0.XI1<7>.XI7<5>.NET_001 XI1.XI0.XI1<7>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_24 XI1.XI0.XI1<7>.XI7<5>.NET_004
+ XI1.XI0.XI1<7>.XI7<5>.NET_000 XI1.XI0.XI1<7>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<5>.NET_005
+ XI1.XI0.XI1<7>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<5>.NET_003
+ XI1.XI0.XI1<7>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_89_4 REG_DATA_7<5> XI1.XI0.XI1<7>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<5>.MM_i_55 XI1.XI0.XI1<7>.XI7<5>.NET_001
+ XI1.XI0.XI1<7>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_61 XI1.XI0.XI1<7>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_66 XI1.XI0.XI1<7>.XI7<5>.NET_003
+ XI1.XI0.XI1<7>.XI7<5>.NET_000 XI1.XI0.XI1<7>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_72 XI1.XI0.XI1<7>.XI7<5>.NET_007
+ XI1.XI0.XI1<7>.XI7<5>.NET_001 XI1.XI0.XI1<7>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<5>.NET_005
+ XI1.XI0.XI1<7>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<5>.NET_003
+ XI1.XI0.XI1<7>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_41_11 REG_DATA_7<4> XI1.XI0.XI1<7>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<4>.MM_i_7 XI1.XI0.XI1<7>.XI7<4>.NET_001
+ XI1.XI0.XI1<7>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_13 XI1.XI0.XI1<7>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_18 XI1.XI0.XI1<7>.XI7<4>.NET_003
+ XI1.XI0.XI1<7>.XI7<4>.NET_001 XI1.XI0.XI1<7>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_24 XI1.XI0.XI1<7>.XI7<4>.NET_004
+ XI1.XI0.XI1<7>.XI7<4>.NET_000 XI1.XI0.XI1<7>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<4>.NET_005
+ XI1.XI0.XI1<7>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<4>.NET_003
+ XI1.XI0.XI1<7>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_89_4 REG_DATA_7<4> XI1.XI0.XI1<7>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<4>.MM_i_55 XI1.XI0.XI1<7>.XI7<4>.NET_001
+ XI1.XI0.XI1<7>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_61 XI1.XI0.XI1<7>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_66 XI1.XI0.XI1<7>.XI7<4>.NET_003
+ XI1.XI0.XI1<7>.XI7<4>.NET_000 XI1.XI0.XI1<7>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_72 XI1.XI0.XI1<7>.XI7<4>.NET_007
+ XI1.XI0.XI1<7>.XI7<4>.NET_001 XI1.XI0.XI1<7>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<4>.NET_005
+ XI1.XI0.XI1<7>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<4>.NET_003
+ XI1.XI0.XI1<7>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_41_11 REG_DATA_7<11> XI1.XI0.XI1<7>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<11>.MM_i_7 XI1.XI0.XI1<7>.XI7<11>.NET_001
+ XI1.XI0.XI1<7>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_13 XI1.XI0.XI1<7>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_18 XI1.XI0.XI1<7>.XI7<11>.NET_003
+ XI1.XI0.XI1<7>.XI7<11>.NET_001 XI1.XI0.XI1<7>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_24 XI1.XI0.XI1<7>.XI7<11>.NET_004
+ XI1.XI0.XI1<7>.XI7<11>.NET_000 XI1.XI0.XI1<7>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<11>.NET_005
+ XI1.XI0.XI1<7>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<11>.NET_003
+ XI1.XI0.XI1<7>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_89_4 REG_DATA_7<11> XI1.XI0.XI1<7>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<11>.MM_i_55 XI1.XI0.XI1<7>.XI7<11>.NET_001
+ XI1.XI0.XI1<7>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_61 XI1.XI0.XI1<7>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_66 XI1.XI0.XI1<7>.XI7<11>.NET_003
+ XI1.XI0.XI1<7>.XI7<11>.NET_000 XI1.XI0.XI1<7>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_72 XI1.XI0.XI1<7>.XI7<11>.NET_007
+ XI1.XI0.XI1<7>.XI7<11>.NET_001 XI1.XI0.XI1<7>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<11>.NET_005
+ XI1.XI0.XI1<7>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<11>.NET_003
+ XI1.XI0.XI1<7>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_41_11 REG_DATA_7<10> XI1.XI0.XI1<7>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<10>.MM_i_7 XI1.XI0.XI1<7>.XI7<10>.NET_001
+ XI1.XI0.XI1<7>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_13 XI1.XI0.XI1<7>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_18 XI1.XI0.XI1<7>.XI7<10>.NET_003
+ XI1.XI0.XI1<7>.XI7<10>.NET_001 XI1.XI0.XI1<7>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_24 XI1.XI0.XI1<7>.XI7<10>.NET_004
+ XI1.XI0.XI1<7>.XI7<10>.NET_000 XI1.XI0.XI1<7>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<10>.NET_005
+ XI1.XI0.XI1<7>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<10>.NET_003
+ XI1.XI0.XI1<7>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_89_4 REG_DATA_7<10> XI1.XI0.XI1<7>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<10>.MM_i_55 XI1.XI0.XI1<7>.XI7<10>.NET_001
+ XI1.XI0.XI1<7>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_61 XI1.XI0.XI1<7>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_66 XI1.XI0.XI1<7>.XI7<10>.NET_003
+ XI1.XI0.XI1<7>.XI7<10>.NET_000 XI1.XI0.XI1<7>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_72 XI1.XI0.XI1<7>.XI7<10>.NET_007
+ XI1.XI0.XI1<7>.XI7<10>.NET_001 XI1.XI0.XI1<7>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<10>.NET_005
+ XI1.XI0.XI1<7>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<10>.NET_003
+ XI1.XI0.XI1<7>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_41_11 REG_DATA_7<9> XI1.XI0.XI1<7>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<9>.MM_i_7 XI1.XI0.XI1<7>.XI7<9>.NET_001
+ XI1.XI0.XI1<7>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_13 XI1.XI0.XI1<7>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_18 XI1.XI0.XI1<7>.XI7<9>.NET_003
+ XI1.XI0.XI1<7>.XI7<9>.NET_001 XI1.XI0.XI1<7>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_24 XI1.XI0.XI1<7>.XI7<9>.NET_004
+ XI1.XI0.XI1<7>.XI7<9>.NET_000 XI1.XI0.XI1<7>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<9>.NET_005
+ XI1.XI0.XI1<7>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<9>.NET_003
+ XI1.XI0.XI1<7>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_89_4 REG_DATA_7<9> XI1.XI0.XI1<7>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<9>.MM_i_55 XI1.XI0.XI1<7>.XI7<9>.NET_001
+ XI1.XI0.XI1<7>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_61 XI1.XI0.XI1<7>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_66 XI1.XI0.XI1<7>.XI7<9>.NET_003
+ XI1.XI0.XI1<7>.XI7<9>.NET_000 XI1.XI0.XI1<7>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_72 XI1.XI0.XI1<7>.XI7<9>.NET_007
+ XI1.XI0.XI1<7>.XI7<9>.NET_001 XI1.XI0.XI1<7>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<9>.NET_005
+ XI1.XI0.XI1<7>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<9>.NET_003
+ XI1.XI0.XI1<7>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_41_11 REG_DATA_7<8> XI1.XI0.XI1<7>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<8>.MM_i_7 XI1.XI0.XI1<7>.XI7<8>.NET_001
+ XI1.XI0.XI1<7>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_13 XI1.XI0.XI1<7>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_18 XI1.XI0.XI1<7>.XI7<8>.NET_003
+ XI1.XI0.XI1<7>.XI7<8>.NET_001 XI1.XI0.XI1<7>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_24 XI1.XI0.XI1<7>.XI7<8>.NET_004
+ XI1.XI0.XI1<7>.XI7<8>.NET_000 XI1.XI0.XI1<7>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<8>.NET_005
+ XI1.XI0.XI1<7>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<8>.NET_003
+ XI1.XI0.XI1<7>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_89_4 REG_DATA_7<8> XI1.XI0.XI1<7>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<8>.MM_i_55 XI1.XI0.XI1<7>.XI7<8>.NET_001
+ XI1.XI0.XI1<7>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_61 XI1.XI0.XI1<7>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_66 XI1.XI0.XI1<7>.XI7<8>.NET_003
+ XI1.XI0.XI1<7>.XI7<8>.NET_000 XI1.XI0.XI1<7>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_72 XI1.XI0.XI1<7>.XI7<8>.NET_007
+ XI1.XI0.XI1<7>.XI7<8>.NET_001 XI1.XI0.XI1<7>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<8>.NET_005
+ XI1.XI0.XI1<7>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<8>.NET_003
+ XI1.XI0.XI1<7>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_41_11 REG_DATA_7<15> XI1.XI0.XI1<7>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<15>.MM_i_7 XI1.XI0.XI1<7>.XI7<15>.NET_001
+ XI1.XI0.XI1<7>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_13 XI1.XI0.XI1<7>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_18 XI1.XI0.XI1<7>.XI7<15>.NET_003
+ XI1.XI0.XI1<7>.XI7<15>.NET_001 XI1.XI0.XI1<7>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_24 XI1.XI0.XI1<7>.XI7<15>.NET_004
+ XI1.XI0.XI1<7>.XI7<15>.NET_000 XI1.XI0.XI1<7>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<15>.NET_005
+ XI1.XI0.XI1<7>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<15>.NET_003
+ XI1.XI0.XI1<7>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_89_4 REG_DATA_7<15> XI1.XI0.XI1<7>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<15>.MM_i_55 XI1.XI0.XI1<7>.XI7<15>.NET_001
+ XI1.XI0.XI1<7>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_61 XI1.XI0.XI1<7>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_66 XI1.XI0.XI1<7>.XI7<15>.NET_003
+ XI1.XI0.XI1<7>.XI7<15>.NET_000 XI1.XI0.XI1<7>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_72 XI1.XI0.XI1<7>.XI7<15>.NET_007
+ XI1.XI0.XI1<7>.XI7<15>.NET_001 XI1.XI0.XI1<7>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<15>.NET_005
+ XI1.XI0.XI1<7>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<15>.NET_003
+ XI1.XI0.XI1<7>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_41_11 REG_DATA_7<14> XI1.XI0.XI1<7>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<14>.MM_i_7 XI1.XI0.XI1<7>.XI7<14>.NET_001
+ XI1.XI0.XI1<7>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_13 XI1.XI0.XI1<7>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_18 XI1.XI0.XI1<7>.XI7<14>.NET_003
+ XI1.XI0.XI1<7>.XI7<14>.NET_001 XI1.XI0.XI1<7>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_24 XI1.XI0.XI1<7>.XI7<14>.NET_004
+ XI1.XI0.XI1<7>.XI7<14>.NET_000 XI1.XI0.XI1<7>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<14>.NET_005
+ XI1.XI0.XI1<7>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<14>.NET_003
+ XI1.XI0.XI1<7>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_89_4 REG_DATA_7<14> XI1.XI0.XI1<7>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<14>.MM_i_55 XI1.XI0.XI1<7>.XI7<14>.NET_001
+ XI1.XI0.XI1<7>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_61 XI1.XI0.XI1<7>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_66 XI1.XI0.XI1<7>.XI7<14>.NET_003
+ XI1.XI0.XI1<7>.XI7<14>.NET_000 XI1.XI0.XI1<7>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_72 XI1.XI0.XI1<7>.XI7<14>.NET_007
+ XI1.XI0.XI1<7>.XI7<14>.NET_001 XI1.XI0.XI1<7>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<14>.NET_005
+ XI1.XI0.XI1<7>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<14>.NET_003
+ XI1.XI0.XI1<7>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_41_11 REG_DATA_7<13> XI1.XI0.XI1<7>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<13>.MM_i_7 XI1.XI0.XI1<7>.XI7<13>.NET_001
+ XI1.XI0.XI1<7>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_13 XI1.XI0.XI1<7>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_18 XI1.XI0.XI1<7>.XI7<13>.NET_003
+ XI1.XI0.XI1<7>.XI7<13>.NET_001 XI1.XI0.XI1<7>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_24 XI1.XI0.XI1<7>.XI7<13>.NET_004
+ XI1.XI0.XI1<7>.XI7<13>.NET_000 XI1.XI0.XI1<7>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<13>.NET_005
+ XI1.XI0.XI1<7>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<13>.NET_003
+ XI1.XI0.XI1<7>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_89_4 REG_DATA_7<13> XI1.XI0.XI1<7>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<13>.MM_i_55 XI1.XI0.XI1<7>.XI7<13>.NET_001
+ XI1.XI0.XI1<7>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_61 XI1.XI0.XI1<7>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_66 XI1.XI0.XI1<7>.XI7<13>.NET_003
+ XI1.XI0.XI1<7>.XI7<13>.NET_000 XI1.XI0.XI1<7>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_72 XI1.XI0.XI1<7>.XI7<13>.NET_007
+ XI1.XI0.XI1<7>.XI7<13>.NET_001 XI1.XI0.XI1<7>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<13>.NET_005
+ XI1.XI0.XI1<7>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<13>.NET_003
+ XI1.XI0.XI1<7>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_41_11 REG_DATA_7<12> XI1.XI0.XI1<7>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<7>.XI7<12>.MM_i_7 XI1.XI0.XI1<7>.XI7<12>.NET_001
+ XI1.XI0.XI1<7>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_13 XI1.XI0.XI1<7>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_18 XI1.XI0.XI1<7>.XI7<12>.NET_003
+ XI1.XI0.XI1<7>.XI7<12>.NET_001 XI1.XI0.XI1<7>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_24 XI1.XI0.XI1<7>.XI7<12>.NET_004
+ XI1.XI0.XI1<7>.XI7<12>.NET_000 XI1.XI0.XI1<7>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<7>.XI7<12>.NET_005
+ XI1.XI0.XI1<7>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<7>.XI7<12>.NET_003
+ XI1.XI0.XI1<7>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<7>
+ XI1.XI0.XI1<7>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_89_4 REG_DATA_7<12> XI1.XI0.XI1<7>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<7>.XI7<12>.MM_i_55 XI1.XI0.XI1<7>.XI7<12>.NET_001
+ XI1.XI0.XI1<7>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_61 XI1.XI0.XI1<7>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_66 XI1.XI0.XI1<7>.XI7<12>.NET_003
+ XI1.XI0.XI1<7>.XI7<12>.NET_000 XI1.XI0.XI1<7>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_72 XI1.XI0.XI1<7>.XI7<12>.NET_007
+ XI1.XI0.XI1<7>.XI7<12>.NET_001 XI1.XI0.XI1<7>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<7>.XI7<12>.NET_005
+ XI1.XI0.XI1<7>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<7>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<7>.XI7<12>.NET_003
+ XI1.XI0.XI1<7>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_41_11 REG_DATA_6<3> XI1.XI0.XI1<6>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<3>.MM_i_7 XI1.XI0.XI1<6>.XI7<3>.NET_001
+ XI1.XI0.XI1<6>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_13 XI1.XI0.XI1<6>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_18 XI1.XI0.XI1<6>.XI7<3>.NET_003
+ XI1.XI0.XI1<6>.XI7<3>.NET_001 XI1.XI0.XI1<6>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_24 XI1.XI0.XI1<6>.XI7<3>.NET_004
+ XI1.XI0.XI1<6>.XI7<3>.NET_000 XI1.XI0.XI1<6>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<3>.NET_005
+ XI1.XI0.XI1<6>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<3>.NET_003
+ XI1.XI0.XI1<6>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_89_4 REG_DATA_6<3> XI1.XI0.XI1<6>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<3>.MM_i_55 XI1.XI0.XI1<6>.XI7<3>.NET_001
+ XI1.XI0.XI1<6>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_61 XI1.XI0.XI1<6>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_66 XI1.XI0.XI1<6>.XI7<3>.NET_003
+ XI1.XI0.XI1<6>.XI7<3>.NET_000 XI1.XI0.XI1<6>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_72 XI1.XI0.XI1<6>.XI7<3>.NET_007
+ XI1.XI0.XI1<6>.XI7<3>.NET_001 XI1.XI0.XI1<6>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<3>.NET_005
+ XI1.XI0.XI1<6>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<3>.NET_003
+ XI1.XI0.XI1<6>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_41_11 REG_DATA_6<2> XI1.XI0.XI1<6>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<2>.MM_i_7 XI1.XI0.XI1<6>.XI7<2>.NET_001
+ XI1.XI0.XI1<6>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_13 XI1.XI0.XI1<6>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_18 XI1.XI0.XI1<6>.XI7<2>.NET_003
+ XI1.XI0.XI1<6>.XI7<2>.NET_001 XI1.XI0.XI1<6>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_24 XI1.XI0.XI1<6>.XI7<2>.NET_004
+ XI1.XI0.XI1<6>.XI7<2>.NET_000 XI1.XI0.XI1<6>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<2>.NET_005
+ XI1.XI0.XI1<6>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<2>.NET_003
+ XI1.XI0.XI1<6>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_89_4 REG_DATA_6<2> XI1.XI0.XI1<6>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<2>.MM_i_55 XI1.XI0.XI1<6>.XI7<2>.NET_001
+ XI1.XI0.XI1<6>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_61 XI1.XI0.XI1<6>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_66 XI1.XI0.XI1<6>.XI7<2>.NET_003
+ XI1.XI0.XI1<6>.XI7<2>.NET_000 XI1.XI0.XI1<6>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_72 XI1.XI0.XI1<6>.XI7<2>.NET_007
+ XI1.XI0.XI1<6>.XI7<2>.NET_001 XI1.XI0.XI1<6>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<2>.NET_005
+ XI1.XI0.XI1<6>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<2>.NET_003
+ XI1.XI0.XI1<6>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_41_11 REG_DATA_6<1> XI1.XI0.XI1<6>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<1>.MM_i_7 XI1.XI0.XI1<6>.XI7<1>.NET_001
+ XI1.XI0.XI1<6>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_13 XI1.XI0.XI1<6>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_18 XI1.XI0.XI1<6>.XI7<1>.NET_003
+ XI1.XI0.XI1<6>.XI7<1>.NET_001 XI1.XI0.XI1<6>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_24 XI1.XI0.XI1<6>.XI7<1>.NET_004
+ XI1.XI0.XI1<6>.XI7<1>.NET_000 XI1.XI0.XI1<6>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<1>.NET_005
+ XI1.XI0.XI1<6>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<1>.NET_003
+ XI1.XI0.XI1<6>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_89_4 REG_DATA_6<1> XI1.XI0.XI1<6>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<1>.MM_i_55 XI1.XI0.XI1<6>.XI7<1>.NET_001
+ XI1.XI0.XI1<6>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_61 XI1.XI0.XI1<6>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_66 XI1.XI0.XI1<6>.XI7<1>.NET_003
+ XI1.XI0.XI1<6>.XI7<1>.NET_000 XI1.XI0.XI1<6>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_72 XI1.XI0.XI1<6>.XI7<1>.NET_007
+ XI1.XI0.XI1<6>.XI7<1>.NET_001 XI1.XI0.XI1<6>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<1>.NET_005
+ XI1.XI0.XI1<6>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<1>.NET_003
+ XI1.XI0.XI1<6>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_41_11 REG_DATA_6<0> XI1.XI0.XI1<6>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<0>.MM_i_7 XI1.XI0.XI1<6>.XI7<0>.NET_001
+ XI1.XI0.XI1<6>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_13 XI1.XI0.XI1<6>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_18 XI1.XI0.XI1<6>.XI7<0>.NET_003
+ XI1.XI0.XI1<6>.XI7<0>.NET_001 XI1.XI0.XI1<6>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_24 XI1.XI0.XI1<6>.XI7<0>.NET_004
+ XI1.XI0.XI1<6>.XI7<0>.NET_000 XI1.XI0.XI1<6>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<0>.NET_005
+ XI1.XI0.XI1<6>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<0>.NET_003
+ XI1.XI0.XI1<6>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_89_4 REG_DATA_6<0> XI1.XI0.XI1<6>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<0>.MM_i_55 XI1.XI0.XI1<6>.XI7<0>.NET_001
+ XI1.XI0.XI1<6>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_61 XI1.XI0.XI1<6>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_66 XI1.XI0.XI1<6>.XI7<0>.NET_003
+ XI1.XI0.XI1<6>.XI7<0>.NET_000 XI1.XI0.XI1<6>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_72 XI1.XI0.XI1<6>.XI7<0>.NET_007
+ XI1.XI0.XI1<6>.XI7<0>.NET_001 XI1.XI0.XI1<6>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<0>.NET_005
+ XI1.XI0.XI1<6>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<0>.NET_003
+ XI1.XI0.XI1<6>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_41_11 REG_DATA_6<7> XI1.XI0.XI1<6>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<7>.MM_i_7 XI1.XI0.XI1<6>.XI7<7>.NET_001
+ XI1.XI0.XI1<6>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_13 XI1.XI0.XI1<6>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_18 XI1.XI0.XI1<6>.XI7<7>.NET_003
+ XI1.XI0.XI1<6>.XI7<7>.NET_001 XI1.XI0.XI1<6>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_24 XI1.XI0.XI1<6>.XI7<7>.NET_004
+ XI1.XI0.XI1<6>.XI7<7>.NET_000 XI1.XI0.XI1<6>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<7>.NET_005
+ XI1.XI0.XI1<6>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<7>.NET_003
+ XI1.XI0.XI1<6>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_89_4 REG_DATA_6<7> XI1.XI0.XI1<6>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<7>.MM_i_55 XI1.XI0.XI1<6>.XI7<7>.NET_001
+ XI1.XI0.XI1<6>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_61 XI1.XI0.XI1<6>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_66 XI1.XI0.XI1<6>.XI7<7>.NET_003
+ XI1.XI0.XI1<6>.XI7<7>.NET_000 XI1.XI0.XI1<6>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_72 XI1.XI0.XI1<6>.XI7<7>.NET_007
+ XI1.XI0.XI1<6>.XI7<7>.NET_001 XI1.XI0.XI1<6>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<7>.NET_005
+ XI1.XI0.XI1<6>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<7>.NET_003
+ XI1.XI0.XI1<6>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_41_11 REG_DATA_6<6> XI1.XI0.XI1<6>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<6>.MM_i_7 XI1.XI0.XI1<6>.XI7<6>.NET_001
+ XI1.XI0.XI1<6>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_13 XI1.XI0.XI1<6>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_18 XI1.XI0.XI1<6>.XI7<6>.NET_003
+ XI1.XI0.XI1<6>.XI7<6>.NET_001 XI1.XI0.XI1<6>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_24 XI1.XI0.XI1<6>.XI7<6>.NET_004
+ XI1.XI0.XI1<6>.XI7<6>.NET_000 XI1.XI0.XI1<6>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<6>.NET_005
+ XI1.XI0.XI1<6>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<6>.NET_003
+ XI1.XI0.XI1<6>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_89_4 REG_DATA_6<6> XI1.XI0.XI1<6>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<6>.MM_i_55 XI1.XI0.XI1<6>.XI7<6>.NET_001
+ XI1.XI0.XI1<6>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_61 XI1.XI0.XI1<6>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_66 XI1.XI0.XI1<6>.XI7<6>.NET_003
+ XI1.XI0.XI1<6>.XI7<6>.NET_000 XI1.XI0.XI1<6>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_72 XI1.XI0.XI1<6>.XI7<6>.NET_007
+ XI1.XI0.XI1<6>.XI7<6>.NET_001 XI1.XI0.XI1<6>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<6>.NET_005
+ XI1.XI0.XI1<6>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<6>.NET_003
+ XI1.XI0.XI1<6>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_41_11 REG_DATA_6<5> XI1.XI0.XI1<6>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<5>.MM_i_7 XI1.XI0.XI1<6>.XI7<5>.NET_001
+ XI1.XI0.XI1<6>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_13 XI1.XI0.XI1<6>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_18 XI1.XI0.XI1<6>.XI7<5>.NET_003
+ XI1.XI0.XI1<6>.XI7<5>.NET_001 XI1.XI0.XI1<6>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_24 XI1.XI0.XI1<6>.XI7<5>.NET_004
+ XI1.XI0.XI1<6>.XI7<5>.NET_000 XI1.XI0.XI1<6>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<5>.NET_005
+ XI1.XI0.XI1<6>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<5>.NET_003
+ XI1.XI0.XI1<6>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_89_4 REG_DATA_6<5> XI1.XI0.XI1<6>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<5>.MM_i_55 XI1.XI0.XI1<6>.XI7<5>.NET_001
+ XI1.XI0.XI1<6>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_61 XI1.XI0.XI1<6>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_66 XI1.XI0.XI1<6>.XI7<5>.NET_003
+ XI1.XI0.XI1<6>.XI7<5>.NET_000 XI1.XI0.XI1<6>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_72 XI1.XI0.XI1<6>.XI7<5>.NET_007
+ XI1.XI0.XI1<6>.XI7<5>.NET_001 XI1.XI0.XI1<6>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<5>.NET_005
+ XI1.XI0.XI1<6>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<5>.NET_003
+ XI1.XI0.XI1<6>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_41_11 REG_DATA_6<4> XI1.XI0.XI1<6>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<4>.MM_i_7 XI1.XI0.XI1<6>.XI7<4>.NET_001
+ XI1.XI0.XI1<6>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_13 XI1.XI0.XI1<6>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_18 XI1.XI0.XI1<6>.XI7<4>.NET_003
+ XI1.XI0.XI1<6>.XI7<4>.NET_001 XI1.XI0.XI1<6>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_24 XI1.XI0.XI1<6>.XI7<4>.NET_004
+ XI1.XI0.XI1<6>.XI7<4>.NET_000 XI1.XI0.XI1<6>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<4>.NET_005
+ XI1.XI0.XI1<6>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<4>.NET_003
+ XI1.XI0.XI1<6>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_89_4 REG_DATA_6<4> XI1.XI0.XI1<6>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<4>.MM_i_55 XI1.XI0.XI1<6>.XI7<4>.NET_001
+ XI1.XI0.XI1<6>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_61 XI1.XI0.XI1<6>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_66 XI1.XI0.XI1<6>.XI7<4>.NET_003
+ XI1.XI0.XI1<6>.XI7<4>.NET_000 XI1.XI0.XI1<6>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_72 XI1.XI0.XI1<6>.XI7<4>.NET_007
+ XI1.XI0.XI1<6>.XI7<4>.NET_001 XI1.XI0.XI1<6>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<4>.NET_005
+ XI1.XI0.XI1<6>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<4>.NET_003
+ XI1.XI0.XI1<6>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_41_11 REG_DATA_6<11> XI1.XI0.XI1<6>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<11>.MM_i_7 XI1.XI0.XI1<6>.XI7<11>.NET_001
+ XI1.XI0.XI1<6>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_13 XI1.XI0.XI1<6>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_18 XI1.XI0.XI1<6>.XI7<11>.NET_003
+ XI1.XI0.XI1<6>.XI7<11>.NET_001 XI1.XI0.XI1<6>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_24 XI1.XI0.XI1<6>.XI7<11>.NET_004
+ XI1.XI0.XI1<6>.XI7<11>.NET_000 XI1.XI0.XI1<6>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<11>.NET_005
+ XI1.XI0.XI1<6>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<11>.NET_003
+ XI1.XI0.XI1<6>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_89_4 REG_DATA_6<11> XI1.XI0.XI1<6>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<11>.MM_i_55 XI1.XI0.XI1<6>.XI7<11>.NET_001
+ XI1.XI0.XI1<6>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_61 XI1.XI0.XI1<6>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_66 XI1.XI0.XI1<6>.XI7<11>.NET_003
+ XI1.XI0.XI1<6>.XI7<11>.NET_000 XI1.XI0.XI1<6>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_72 XI1.XI0.XI1<6>.XI7<11>.NET_007
+ XI1.XI0.XI1<6>.XI7<11>.NET_001 XI1.XI0.XI1<6>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<11>.NET_005
+ XI1.XI0.XI1<6>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<11>.NET_003
+ XI1.XI0.XI1<6>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_41_11 REG_DATA_6<10> XI1.XI0.XI1<6>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<10>.MM_i_7 XI1.XI0.XI1<6>.XI7<10>.NET_001
+ XI1.XI0.XI1<6>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_13 XI1.XI0.XI1<6>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_18 XI1.XI0.XI1<6>.XI7<10>.NET_003
+ XI1.XI0.XI1<6>.XI7<10>.NET_001 XI1.XI0.XI1<6>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_24 XI1.XI0.XI1<6>.XI7<10>.NET_004
+ XI1.XI0.XI1<6>.XI7<10>.NET_000 XI1.XI0.XI1<6>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<10>.NET_005
+ XI1.XI0.XI1<6>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<10>.NET_003
+ XI1.XI0.XI1<6>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_89_4 REG_DATA_6<10> XI1.XI0.XI1<6>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<10>.MM_i_55 XI1.XI0.XI1<6>.XI7<10>.NET_001
+ XI1.XI0.XI1<6>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_61 XI1.XI0.XI1<6>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_66 XI1.XI0.XI1<6>.XI7<10>.NET_003
+ XI1.XI0.XI1<6>.XI7<10>.NET_000 XI1.XI0.XI1<6>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_72 XI1.XI0.XI1<6>.XI7<10>.NET_007
+ XI1.XI0.XI1<6>.XI7<10>.NET_001 XI1.XI0.XI1<6>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<10>.NET_005
+ XI1.XI0.XI1<6>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<10>.NET_003
+ XI1.XI0.XI1<6>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_41_11 REG_DATA_6<9> XI1.XI0.XI1<6>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<9>.MM_i_7 XI1.XI0.XI1<6>.XI7<9>.NET_001
+ XI1.XI0.XI1<6>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_13 XI1.XI0.XI1<6>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_18 XI1.XI0.XI1<6>.XI7<9>.NET_003
+ XI1.XI0.XI1<6>.XI7<9>.NET_001 XI1.XI0.XI1<6>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_24 XI1.XI0.XI1<6>.XI7<9>.NET_004
+ XI1.XI0.XI1<6>.XI7<9>.NET_000 XI1.XI0.XI1<6>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<9>.NET_005
+ XI1.XI0.XI1<6>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<9>.NET_003
+ XI1.XI0.XI1<6>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_89_4 REG_DATA_6<9> XI1.XI0.XI1<6>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<9>.MM_i_55 XI1.XI0.XI1<6>.XI7<9>.NET_001
+ XI1.XI0.XI1<6>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_61 XI1.XI0.XI1<6>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_66 XI1.XI0.XI1<6>.XI7<9>.NET_003
+ XI1.XI0.XI1<6>.XI7<9>.NET_000 XI1.XI0.XI1<6>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_72 XI1.XI0.XI1<6>.XI7<9>.NET_007
+ XI1.XI0.XI1<6>.XI7<9>.NET_001 XI1.XI0.XI1<6>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<9>.NET_005
+ XI1.XI0.XI1<6>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<9>.NET_003
+ XI1.XI0.XI1<6>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_41_11 REG_DATA_6<8> XI1.XI0.XI1<6>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<8>.MM_i_7 XI1.XI0.XI1<6>.XI7<8>.NET_001
+ XI1.XI0.XI1<6>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_13 XI1.XI0.XI1<6>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_18 XI1.XI0.XI1<6>.XI7<8>.NET_003
+ XI1.XI0.XI1<6>.XI7<8>.NET_001 XI1.XI0.XI1<6>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_24 XI1.XI0.XI1<6>.XI7<8>.NET_004
+ XI1.XI0.XI1<6>.XI7<8>.NET_000 XI1.XI0.XI1<6>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<8>.NET_005
+ XI1.XI0.XI1<6>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<8>.NET_003
+ XI1.XI0.XI1<6>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_89_4 REG_DATA_6<8> XI1.XI0.XI1<6>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<8>.MM_i_55 XI1.XI0.XI1<6>.XI7<8>.NET_001
+ XI1.XI0.XI1<6>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_61 XI1.XI0.XI1<6>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_66 XI1.XI0.XI1<6>.XI7<8>.NET_003
+ XI1.XI0.XI1<6>.XI7<8>.NET_000 XI1.XI0.XI1<6>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_72 XI1.XI0.XI1<6>.XI7<8>.NET_007
+ XI1.XI0.XI1<6>.XI7<8>.NET_001 XI1.XI0.XI1<6>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<8>.NET_005
+ XI1.XI0.XI1<6>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<8>.NET_003
+ XI1.XI0.XI1<6>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_41_11 REG_DATA_6<15> XI1.XI0.XI1<6>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<15>.MM_i_7 XI1.XI0.XI1<6>.XI7<15>.NET_001
+ XI1.XI0.XI1<6>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_13 XI1.XI0.XI1<6>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_18 XI1.XI0.XI1<6>.XI7<15>.NET_003
+ XI1.XI0.XI1<6>.XI7<15>.NET_001 XI1.XI0.XI1<6>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_24 XI1.XI0.XI1<6>.XI7<15>.NET_004
+ XI1.XI0.XI1<6>.XI7<15>.NET_000 XI1.XI0.XI1<6>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<15>.NET_005
+ XI1.XI0.XI1<6>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<15>.NET_003
+ XI1.XI0.XI1<6>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_89_4 REG_DATA_6<15> XI1.XI0.XI1<6>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<15>.MM_i_55 XI1.XI0.XI1<6>.XI7<15>.NET_001
+ XI1.XI0.XI1<6>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_61 XI1.XI0.XI1<6>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_66 XI1.XI0.XI1<6>.XI7<15>.NET_003
+ XI1.XI0.XI1<6>.XI7<15>.NET_000 XI1.XI0.XI1<6>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_72 XI1.XI0.XI1<6>.XI7<15>.NET_007
+ XI1.XI0.XI1<6>.XI7<15>.NET_001 XI1.XI0.XI1<6>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<15>.NET_005
+ XI1.XI0.XI1<6>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<15>.NET_003
+ XI1.XI0.XI1<6>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_41_11 REG_DATA_6<14> XI1.XI0.XI1<6>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<14>.MM_i_7 XI1.XI0.XI1<6>.XI7<14>.NET_001
+ XI1.XI0.XI1<6>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_13 XI1.XI0.XI1<6>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_18 XI1.XI0.XI1<6>.XI7<14>.NET_003
+ XI1.XI0.XI1<6>.XI7<14>.NET_001 XI1.XI0.XI1<6>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_24 XI1.XI0.XI1<6>.XI7<14>.NET_004
+ XI1.XI0.XI1<6>.XI7<14>.NET_000 XI1.XI0.XI1<6>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<14>.NET_005
+ XI1.XI0.XI1<6>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<14>.NET_003
+ XI1.XI0.XI1<6>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_89_4 REG_DATA_6<14> XI1.XI0.XI1<6>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<14>.MM_i_55 XI1.XI0.XI1<6>.XI7<14>.NET_001
+ XI1.XI0.XI1<6>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_61 XI1.XI0.XI1<6>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_66 XI1.XI0.XI1<6>.XI7<14>.NET_003
+ XI1.XI0.XI1<6>.XI7<14>.NET_000 XI1.XI0.XI1<6>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_72 XI1.XI0.XI1<6>.XI7<14>.NET_007
+ XI1.XI0.XI1<6>.XI7<14>.NET_001 XI1.XI0.XI1<6>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<14>.NET_005
+ XI1.XI0.XI1<6>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<14>.NET_003
+ XI1.XI0.XI1<6>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_41_11 REG_DATA_6<13> XI1.XI0.XI1<6>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<13>.MM_i_7 XI1.XI0.XI1<6>.XI7<13>.NET_001
+ XI1.XI0.XI1<6>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_13 XI1.XI0.XI1<6>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_18 XI1.XI0.XI1<6>.XI7<13>.NET_003
+ XI1.XI0.XI1<6>.XI7<13>.NET_001 XI1.XI0.XI1<6>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_24 XI1.XI0.XI1<6>.XI7<13>.NET_004
+ XI1.XI0.XI1<6>.XI7<13>.NET_000 XI1.XI0.XI1<6>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<13>.NET_005
+ XI1.XI0.XI1<6>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<13>.NET_003
+ XI1.XI0.XI1<6>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_89_4 REG_DATA_6<13> XI1.XI0.XI1<6>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<13>.MM_i_55 XI1.XI0.XI1<6>.XI7<13>.NET_001
+ XI1.XI0.XI1<6>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_61 XI1.XI0.XI1<6>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_66 XI1.XI0.XI1<6>.XI7<13>.NET_003
+ XI1.XI0.XI1<6>.XI7<13>.NET_000 XI1.XI0.XI1<6>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_72 XI1.XI0.XI1<6>.XI7<13>.NET_007
+ XI1.XI0.XI1<6>.XI7<13>.NET_001 XI1.XI0.XI1<6>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<13>.NET_005
+ XI1.XI0.XI1<6>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<13>.NET_003
+ XI1.XI0.XI1<6>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_41_11 REG_DATA_6<12> XI1.XI0.XI1<6>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<6>.XI7<12>.MM_i_7 XI1.XI0.XI1<6>.XI7<12>.NET_001
+ XI1.XI0.XI1<6>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_13 XI1.XI0.XI1<6>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_18 XI1.XI0.XI1<6>.XI7<12>.NET_003
+ XI1.XI0.XI1<6>.XI7<12>.NET_001 XI1.XI0.XI1<6>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_24 XI1.XI0.XI1<6>.XI7<12>.NET_004
+ XI1.XI0.XI1<6>.XI7<12>.NET_000 XI1.XI0.XI1<6>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<6>.XI7<12>.NET_005
+ XI1.XI0.XI1<6>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<6>.XI7<12>.NET_003
+ XI1.XI0.XI1<6>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<6>
+ XI1.XI0.XI1<6>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_89_4 REG_DATA_6<12> XI1.XI0.XI1<6>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<6>.XI7<12>.MM_i_55 XI1.XI0.XI1<6>.XI7<12>.NET_001
+ XI1.XI0.XI1<6>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_61 XI1.XI0.XI1<6>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_66 XI1.XI0.XI1<6>.XI7<12>.NET_003
+ XI1.XI0.XI1<6>.XI7<12>.NET_000 XI1.XI0.XI1<6>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_72 XI1.XI0.XI1<6>.XI7<12>.NET_007
+ XI1.XI0.XI1<6>.XI7<12>.NET_001 XI1.XI0.XI1<6>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<6>.XI7<12>.NET_005
+ XI1.XI0.XI1<6>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<6>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<6>.XI7<12>.NET_003
+ XI1.XI0.XI1<6>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_41_11 REG_DATA_5<3> XI1.XI0.XI1<5>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<3>.MM_i_7 XI1.XI0.XI1<5>.XI7<3>.NET_001
+ XI1.XI0.XI1<5>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_13 XI1.XI0.XI1<5>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_18 XI1.XI0.XI1<5>.XI7<3>.NET_003
+ XI1.XI0.XI1<5>.XI7<3>.NET_001 XI1.XI0.XI1<5>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_24 XI1.XI0.XI1<5>.XI7<3>.NET_004
+ XI1.XI0.XI1<5>.XI7<3>.NET_000 XI1.XI0.XI1<5>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<3>.NET_005
+ XI1.XI0.XI1<5>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<3>.NET_003
+ XI1.XI0.XI1<5>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_89_4 REG_DATA_5<3> XI1.XI0.XI1<5>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<3>.MM_i_55 XI1.XI0.XI1<5>.XI7<3>.NET_001
+ XI1.XI0.XI1<5>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_61 XI1.XI0.XI1<5>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_66 XI1.XI0.XI1<5>.XI7<3>.NET_003
+ XI1.XI0.XI1<5>.XI7<3>.NET_000 XI1.XI0.XI1<5>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_72 XI1.XI0.XI1<5>.XI7<3>.NET_007
+ XI1.XI0.XI1<5>.XI7<3>.NET_001 XI1.XI0.XI1<5>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<3>.NET_005
+ XI1.XI0.XI1<5>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<3>.NET_003
+ XI1.XI0.XI1<5>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_41_11 REG_DATA_5<2> XI1.XI0.XI1<5>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<2>.MM_i_7 XI1.XI0.XI1<5>.XI7<2>.NET_001
+ XI1.XI0.XI1<5>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_13 XI1.XI0.XI1<5>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_18 XI1.XI0.XI1<5>.XI7<2>.NET_003
+ XI1.XI0.XI1<5>.XI7<2>.NET_001 XI1.XI0.XI1<5>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_24 XI1.XI0.XI1<5>.XI7<2>.NET_004
+ XI1.XI0.XI1<5>.XI7<2>.NET_000 XI1.XI0.XI1<5>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<2>.NET_005
+ XI1.XI0.XI1<5>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<2>.NET_003
+ XI1.XI0.XI1<5>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_89_4 REG_DATA_5<2> XI1.XI0.XI1<5>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<2>.MM_i_55 XI1.XI0.XI1<5>.XI7<2>.NET_001
+ XI1.XI0.XI1<5>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_61 XI1.XI0.XI1<5>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_66 XI1.XI0.XI1<5>.XI7<2>.NET_003
+ XI1.XI0.XI1<5>.XI7<2>.NET_000 XI1.XI0.XI1<5>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_72 XI1.XI0.XI1<5>.XI7<2>.NET_007
+ XI1.XI0.XI1<5>.XI7<2>.NET_001 XI1.XI0.XI1<5>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<2>.NET_005
+ XI1.XI0.XI1<5>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<2>.NET_003
+ XI1.XI0.XI1<5>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_41_11 REG_DATA_5<1> XI1.XI0.XI1<5>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<1>.MM_i_7 XI1.XI0.XI1<5>.XI7<1>.NET_001
+ XI1.XI0.XI1<5>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_13 XI1.XI0.XI1<5>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_18 XI1.XI0.XI1<5>.XI7<1>.NET_003
+ XI1.XI0.XI1<5>.XI7<1>.NET_001 XI1.XI0.XI1<5>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_24 XI1.XI0.XI1<5>.XI7<1>.NET_004
+ XI1.XI0.XI1<5>.XI7<1>.NET_000 XI1.XI0.XI1<5>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<1>.NET_005
+ XI1.XI0.XI1<5>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<1>.NET_003
+ XI1.XI0.XI1<5>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_89_4 REG_DATA_5<1> XI1.XI0.XI1<5>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<1>.MM_i_55 XI1.XI0.XI1<5>.XI7<1>.NET_001
+ XI1.XI0.XI1<5>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_61 XI1.XI0.XI1<5>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_66 XI1.XI0.XI1<5>.XI7<1>.NET_003
+ XI1.XI0.XI1<5>.XI7<1>.NET_000 XI1.XI0.XI1<5>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_72 XI1.XI0.XI1<5>.XI7<1>.NET_007
+ XI1.XI0.XI1<5>.XI7<1>.NET_001 XI1.XI0.XI1<5>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<1>.NET_005
+ XI1.XI0.XI1<5>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<1>.NET_003
+ XI1.XI0.XI1<5>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_41_11 REG_DATA_5<0> XI1.XI0.XI1<5>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<0>.MM_i_7 XI1.XI0.XI1<5>.XI7<0>.NET_001
+ XI1.XI0.XI1<5>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_13 XI1.XI0.XI1<5>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_18 XI1.XI0.XI1<5>.XI7<0>.NET_003
+ XI1.XI0.XI1<5>.XI7<0>.NET_001 XI1.XI0.XI1<5>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_24 XI1.XI0.XI1<5>.XI7<0>.NET_004
+ XI1.XI0.XI1<5>.XI7<0>.NET_000 XI1.XI0.XI1<5>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<0>.NET_005
+ XI1.XI0.XI1<5>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<0>.NET_003
+ XI1.XI0.XI1<5>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_89_4 REG_DATA_5<0> XI1.XI0.XI1<5>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<0>.MM_i_55 XI1.XI0.XI1<5>.XI7<0>.NET_001
+ XI1.XI0.XI1<5>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_61 XI1.XI0.XI1<5>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_66 XI1.XI0.XI1<5>.XI7<0>.NET_003
+ XI1.XI0.XI1<5>.XI7<0>.NET_000 XI1.XI0.XI1<5>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_72 XI1.XI0.XI1<5>.XI7<0>.NET_007
+ XI1.XI0.XI1<5>.XI7<0>.NET_001 XI1.XI0.XI1<5>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<0>.NET_005
+ XI1.XI0.XI1<5>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<0>.NET_003
+ XI1.XI0.XI1<5>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_41_11 REG_DATA_5<7> XI1.XI0.XI1<5>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<7>.MM_i_7 XI1.XI0.XI1<5>.XI7<7>.NET_001
+ XI1.XI0.XI1<5>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_13 XI1.XI0.XI1<5>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_18 XI1.XI0.XI1<5>.XI7<7>.NET_003
+ XI1.XI0.XI1<5>.XI7<7>.NET_001 XI1.XI0.XI1<5>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_24 XI1.XI0.XI1<5>.XI7<7>.NET_004
+ XI1.XI0.XI1<5>.XI7<7>.NET_000 XI1.XI0.XI1<5>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<7>.NET_005
+ XI1.XI0.XI1<5>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<7>.NET_003
+ XI1.XI0.XI1<5>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_89_4 REG_DATA_5<7> XI1.XI0.XI1<5>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<7>.MM_i_55 XI1.XI0.XI1<5>.XI7<7>.NET_001
+ XI1.XI0.XI1<5>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_61 XI1.XI0.XI1<5>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_66 XI1.XI0.XI1<5>.XI7<7>.NET_003
+ XI1.XI0.XI1<5>.XI7<7>.NET_000 XI1.XI0.XI1<5>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_72 XI1.XI0.XI1<5>.XI7<7>.NET_007
+ XI1.XI0.XI1<5>.XI7<7>.NET_001 XI1.XI0.XI1<5>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<7>.NET_005
+ XI1.XI0.XI1<5>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<7>.NET_003
+ XI1.XI0.XI1<5>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_41_11 REG_DATA_5<6> XI1.XI0.XI1<5>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<6>.MM_i_7 XI1.XI0.XI1<5>.XI7<6>.NET_001
+ XI1.XI0.XI1<5>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_13 XI1.XI0.XI1<5>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_18 XI1.XI0.XI1<5>.XI7<6>.NET_003
+ XI1.XI0.XI1<5>.XI7<6>.NET_001 XI1.XI0.XI1<5>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_24 XI1.XI0.XI1<5>.XI7<6>.NET_004
+ XI1.XI0.XI1<5>.XI7<6>.NET_000 XI1.XI0.XI1<5>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<6>.NET_005
+ XI1.XI0.XI1<5>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<6>.NET_003
+ XI1.XI0.XI1<5>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_89_4 REG_DATA_5<6> XI1.XI0.XI1<5>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<6>.MM_i_55 XI1.XI0.XI1<5>.XI7<6>.NET_001
+ XI1.XI0.XI1<5>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_61 XI1.XI0.XI1<5>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_66 XI1.XI0.XI1<5>.XI7<6>.NET_003
+ XI1.XI0.XI1<5>.XI7<6>.NET_000 XI1.XI0.XI1<5>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_72 XI1.XI0.XI1<5>.XI7<6>.NET_007
+ XI1.XI0.XI1<5>.XI7<6>.NET_001 XI1.XI0.XI1<5>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<6>.NET_005
+ XI1.XI0.XI1<5>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<6>.NET_003
+ XI1.XI0.XI1<5>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_41_11 REG_DATA_5<5> XI1.XI0.XI1<5>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<5>.MM_i_7 XI1.XI0.XI1<5>.XI7<5>.NET_001
+ XI1.XI0.XI1<5>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_13 XI1.XI0.XI1<5>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_18 XI1.XI0.XI1<5>.XI7<5>.NET_003
+ XI1.XI0.XI1<5>.XI7<5>.NET_001 XI1.XI0.XI1<5>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_24 XI1.XI0.XI1<5>.XI7<5>.NET_004
+ XI1.XI0.XI1<5>.XI7<5>.NET_000 XI1.XI0.XI1<5>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<5>.NET_005
+ XI1.XI0.XI1<5>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<5>.NET_003
+ XI1.XI0.XI1<5>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_89_4 REG_DATA_5<5> XI1.XI0.XI1<5>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<5>.MM_i_55 XI1.XI0.XI1<5>.XI7<5>.NET_001
+ XI1.XI0.XI1<5>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_61 XI1.XI0.XI1<5>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_66 XI1.XI0.XI1<5>.XI7<5>.NET_003
+ XI1.XI0.XI1<5>.XI7<5>.NET_000 XI1.XI0.XI1<5>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_72 XI1.XI0.XI1<5>.XI7<5>.NET_007
+ XI1.XI0.XI1<5>.XI7<5>.NET_001 XI1.XI0.XI1<5>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<5>.NET_005
+ XI1.XI0.XI1<5>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<5>.NET_003
+ XI1.XI0.XI1<5>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_41_11 REG_DATA_5<4> XI1.XI0.XI1<5>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<4>.MM_i_7 XI1.XI0.XI1<5>.XI7<4>.NET_001
+ XI1.XI0.XI1<5>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_13 XI1.XI0.XI1<5>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_18 XI1.XI0.XI1<5>.XI7<4>.NET_003
+ XI1.XI0.XI1<5>.XI7<4>.NET_001 XI1.XI0.XI1<5>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_24 XI1.XI0.XI1<5>.XI7<4>.NET_004
+ XI1.XI0.XI1<5>.XI7<4>.NET_000 XI1.XI0.XI1<5>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<4>.NET_005
+ XI1.XI0.XI1<5>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<4>.NET_003
+ XI1.XI0.XI1<5>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_89_4 REG_DATA_5<4> XI1.XI0.XI1<5>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<4>.MM_i_55 XI1.XI0.XI1<5>.XI7<4>.NET_001
+ XI1.XI0.XI1<5>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_61 XI1.XI0.XI1<5>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_66 XI1.XI0.XI1<5>.XI7<4>.NET_003
+ XI1.XI0.XI1<5>.XI7<4>.NET_000 XI1.XI0.XI1<5>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_72 XI1.XI0.XI1<5>.XI7<4>.NET_007
+ XI1.XI0.XI1<5>.XI7<4>.NET_001 XI1.XI0.XI1<5>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<4>.NET_005
+ XI1.XI0.XI1<5>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<4>.NET_003
+ XI1.XI0.XI1<5>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_41_11 REG_DATA_5<11> XI1.XI0.XI1<5>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<11>.MM_i_7 XI1.XI0.XI1<5>.XI7<11>.NET_001
+ XI1.XI0.XI1<5>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_13 XI1.XI0.XI1<5>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_18 XI1.XI0.XI1<5>.XI7<11>.NET_003
+ XI1.XI0.XI1<5>.XI7<11>.NET_001 XI1.XI0.XI1<5>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_24 XI1.XI0.XI1<5>.XI7<11>.NET_004
+ XI1.XI0.XI1<5>.XI7<11>.NET_000 XI1.XI0.XI1<5>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<11>.NET_005
+ XI1.XI0.XI1<5>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<11>.NET_003
+ XI1.XI0.XI1<5>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_89_4 REG_DATA_5<11> XI1.XI0.XI1<5>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<11>.MM_i_55 XI1.XI0.XI1<5>.XI7<11>.NET_001
+ XI1.XI0.XI1<5>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_61 XI1.XI0.XI1<5>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_66 XI1.XI0.XI1<5>.XI7<11>.NET_003
+ XI1.XI0.XI1<5>.XI7<11>.NET_000 XI1.XI0.XI1<5>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_72 XI1.XI0.XI1<5>.XI7<11>.NET_007
+ XI1.XI0.XI1<5>.XI7<11>.NET_001 XI1.XI0.XI1<5>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<11>.NET_005
+ XI1.XI0.XI1<5>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<11>.NET_003
+ XI1.XI0.XI1<5>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_41_11 REG_DATA_5<10> XI1.XI0.XI1<5>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<10>.MM_i_7 XI1.XI0.XI1<5>.XI7<10>.NET_001
+ XI1.XI0.XI1<5>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_13 XI1.XI0.XI1<5>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_18 XI1.XI0.XI1<5>.XI7<10>.NET_003
+ XI1.XI0.XI1<5>.XI7<10>.NET_001 XI1.XI0.XI1<5>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_24 XI1.XI0.XI1<5>.XI7<10>.NET_004
+ XI1.XI0.XI1<5>.XI7<10>.NET_000 XI1.XI0.XI1<5>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<10>.NET_005
+ XI1.XI0.XI1<5>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<10>.NET_003
+ XI1.XI0.XI1<5>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_89_4 REG_DATA_5<10> XI1.XI0.XI1<5>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<10>.MM_i_55 XI1.XI0.XI1<5>.XI7<10>.NET_001
+ XI1.XI0.XI1<5>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_61 XI1.XI0.XI1<5>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_66 XI1.XI0.XI1<5>.XI7<10>.NET_003
+ XI1.XI0.XI1<5>.XI7<10>.NET_000 XI1.XI0.XI1<5>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_72 XI1.XI0.XI1<5>.XI7<10>.NET_007
+ XI1.XI0.XI1<5>.XI7<10>.NET_001 XI1.XI0.XI1<5>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<10>.NET_005
+ XI1.XI0.XI1<5>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<10>.NET_003
+ XI1.XI0.XI1<5>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_41_11 REG_DATA_5<9> XI1.XI0.XI1<5>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<9>.MM_i_7 XI1.XI0.XI1<5>.XI7<9>.NET_001
+ XI1.XI0.XI1<5>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_13 XI1.XI0.XI1<5>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_18 XI1.XI0.XI1<5>.XI7<9>.NET_003
+ XI1.XI0.XI1<5>.XI7<9>.NET_001 XI1.XI0.XI1<5>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_24 XI1.XI0.XI1<5>.XI7<9>.NET_004
+ XI1.XI0.XI1<5>.XI7<9>.NET_000 XI1.XI0.XI1<5>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<9>.NET_005
+ XI1.XI0.XI1<5>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<9>.NET_003
+ XI1.XI0.XI1<5>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_89_4 REG_DATA_5<9> XI1.XI0.XI1<5>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<9>.MM_i_55 XI1.XI0.XI1<5>.XI7<9>.NET_001
+ XI1.XI0.XI1<5>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_61 XI1.XI0.XI1<5>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_66 XI1.XI0.XI1<5>.XI7<9>.NET_003
+ XI1.XI0.XI1<5>.XI7<9>.NET_000 XI1.XI0.XI1<5>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_72 XI1.XI0.XI1<5>.XI7<9>.NET_007
+ XI1.XI0.XI1<5>.XI7<9>.NET_001 XI1.XI0.XI1<5>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<9>.NET_005
+ XI1.XI0.XI1<5>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<9>.NET_003
+ XI1.XI0.XI1<5>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_41_11 REG_DATA_5<8> XI1.XI0.XI1<5>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<8>.MM_i_7 XI1.XI0.XI1<5>.XI7<8>.NET_001
+ XI1.XI0.XI1<5>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_13 XI1.XI0.XI1<5>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_18 XI1.XI0.XI1<5>.XI7<8>.NET_003
+ XI1.XI0.XI1<5>.XI7<8>.NET_001 XI1.XI0.XI1<5>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_24 XI1.XI0.XI1<5>.XI7<8>.NET_004
+ XI1.XI0.XI1<5>.XI7<8>.NET_000 XI1.XI0.XI1<5>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<8>.NET_005
+ XI1.XI0.XI1<5>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<8>.NET_003
+ XI1.XI0.XI1<5>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_89_4 REG_DATA_5<8> XI1.XI0.XI1<5>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<8>.MM_i_55 XI1.XI0.XI1<5>.XI7<8>.NET_001
+ XI1.XI0.XI1<5>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_61 XI1.XI0.XI1<5>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_66 XI1.XI0.XI1<5>.XI7<8>.NET_003
+ XI1.XI0.XI1<5>.XI7<8>.NET_000 XI1.XI0.XI1<5>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_72 XI1.XI0.XI1<5>.XI7<8>.NET_007
+ XI1.XI0.XI1<5>.XI7<8>.NET_001 XI1.XI0.XI1<5>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<8>.NET_005
+ XI1.XI0.XI1<5>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<8>.NET_003
+ XI1.XI0.XI1<5>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_41_11 REG_DATA_5<15> XI1.XI0.XI1<5>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<15>.MM_i_7 XI1.XI0.XI1<5>.XI7<15>.NET_001
+ XI1.XI0.XI1<5>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_13 XI1.XI0.XI1<5>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_18 XI1.XI0.XI1<5>.XI7<15>.NET_003
+ XI1.XI0.XI1<5>.XI7<15>.NET_001 XI1.XI0.XI1<5>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_24 XI1.XI0.XI1<5>.XI7<15>.NET_004
+ XI1.XI0.XI1<5>.XI7<15>.NET_000 XI1.XI0.XI1<5>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<15>.NET_005
+ XI1.XI0.XI1<5>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<15>.NET_003
+ XI1.XI0.XI1<5>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_89_4 REG_DATA_5<15> XI1.XI0.XI1<5>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<15>.MM_i_55 XI1.XI0.XI1<5>.XI7<15>.NET_001
+ XI1.XI0.XI1<5>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_61 XI1.XI0.XI1<5>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_66 XI1.XI0.XI1<5>.XI7<15>.NET_003
+ XI1.XI0.XI1<5>.XI7<15>.NET_000 XI1.XI0.XI1<5>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_72 XI1.XI0.XI1<5>.XI7<15>.NET_007
+ XI1.XI0.XI1<5>.XI7<15>.NET_001 XI1.XI0.XI1<5>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<15>.NET_005
+ XI1.XI0.XI1<5>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<15>.NET_003
+ XI1.XI0.XI1<5>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_41_11 REG_DATA_5<14> XI1.XI0.XI1<5>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<14>.MM_i_7 XI1.XI0.XI1<5>.XI7<14>.NET_001
+ XI1.XI0.XI1<5>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_13 XI1.XI0.XI1<5>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_18 XI1.XI0.XI1<5>.XI7<14>.NET_003
+ XI1.XI0.XI1<5>.XI7<14>.NET_001 XI1.XI0.XI1<5>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_24 XI1.XI0.XI1<5>.XI7<14>.NET_004
+ XI1.XI0.XI1<5>.XI7<14>.NET_000 XI1.XI0.XI1<5>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<14>.NET_005
+ XI1.XI0.XI1<5>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<14>.NET_003
+ XI1.XI0.XI1<5>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_89_4 REG_DATA_5<14> XI1.XI0.XI1<5>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<14>.MM_i_55 XI1.XI0.XI1<5>.XI7<14>.NET_001
+ XI1.XI0.XI1<5>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_61 XI1.XI0.XI1<5>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_66 XI1.XI0.XI1<5>.XI7<14>.NET_003
+ XI1.XI0.XI1<5>.XI7<14>.NET_000 XI1.XI0.XI1<5>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_72 XI1.XI0.XI1<5>.XI7<14>.NET_007
+ XI1.XI0.XI1<5>.XI7<14>.NET_001 XI1.XI0.XI1<5>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<14>.NET_005
+ XI1.XI0.XI1<5>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<14>.NET_003
+ XI1.XI0.XI1<5>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_41_11 REG_DATA_5<13> XI1.XI0.XI1<5>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<13>.MM_i_7 XI1.XI0.XI1<5>.XI7<13>.NET_001
+ XI1.XI0.XI1<5>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_13 XI1.XI0.XI1<5>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_18 XI1.XI0.XI1<5>.XI7<13>.NET_003
+ XI1.XI0.XI1<5>.XI7<13>.NET_001 XI1.XI0.XI1<5>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_24 XI1.XI0.XI1<5>.XI7<13>.NET_004
+ XI1.XI0.XI1<5>.XI7<13>.NET_000 XI1.XI0.XI1<5>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<13>.NET_005
+ XI1.XI0.XI1<5>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<13>.NET_003
+ XI1.XI0.XI1<5>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_89_4 REG_DATA_5<13> XI1.XI0.XI1<5>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<13>.MM_i_55 XI1.XI0.XI1<5>.XI7<13>.NET_001
+ XI1.XI0.XI1<5>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_61 XI1.XI0.XI1<5>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_66 XI1.XI0.XI1<5>.XI7<13>.NET_003
+ XI1.XI0.XI1<5>.XI7<13>.NET_000 XI1.XI0.XI1<5>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_72 XI1.XI0.XI1<5>.XI7<13>.NET_007
+ XI1.XI0.XI1<5>.XI7<13>.NET_001 XI1.XI0.XI1<5>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<13>.NET_005
+ XI1.XI0.XI1<5>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<13>.NET_003
+ XI1.XI0.XI1<5>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_41_11 REG_DATA_5<12> XI1.XI0.XI1<5>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<5>.XI7<12>.MM_i_7 XI1.XI0.XI1<5>.XI7<12>.NET_001
+ XI1.XI0.XI1<5>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_13 XI1.XI0.XI1<5>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_18 XI1.XI0.XI1<5>.XI7<12>.NET_003
+ XI1.XI0.XI1<5>.XI7<12>.NET_001 XI1.XI0.XI1<5>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_24 XI1.XI0.XI1<5>.XI7<12>.NET_004
+ XI1.XI0.XI1<5>.XI7<12>.NET_000 XI1.XI0.XI1<5>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<5>.XI7<12>.NET_005
+ XI1.XI0.XI1<5>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<5>.XI7<12>.NET_003
+ XI1.XI0.XI1<5>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<5>
+ XI1.XI0.XI1<5>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_89_4 REG_DATA_5<12> XI1.XI0.XI1<5>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<5>.XI7<12>.MM_i_55 XI1.XI0.XI1<5>.XI7<12>.NET_001
+ XI1.XI0.XI1<5>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_61 XI1.XI0.XI1<5>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_66 XI1.XI0.XI1<5>.XI7<12>.NET_003
+ XI1.XI0.XI1<5>.XI7<12>.NET_000 XI1.XI0.XI1<5>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_72 XI1.XI0.XI1<5>.XI7<12>.NET_007
+ XI1.XI0.XI1<5>.XI7<12>.NET_001 XI1.XI0.XI1<5>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<5>.XI7<12>.NET_005
+ XI1.XI0.XI1<5>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<5>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<5>.XI7<12>.NET_003
+ XI1.XI0.XI1<5>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_41_11 REG_DATA_4<3> XI1.XI0.XI1<4>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<3>.MM_i_7 XI1.XI0.XI1<4>.XI7<3>.NET_001
+ XI1.XI0.XI1<4>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_13 XI1.XI0.XI1<4>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_18 XI1.XI0.XI1<4>.XI7<3>.NET_003
+ XI1.XI0.XI1<4>.XI7<3>.NET_001 XI1.XI0.XI1<4>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_24 XI1.XI0.XI1<4>.XI7<3>.NET_004
+ XI1.XI0.XI1<4>.XI7<3>.NET_000 XI1.XI0.XI1<4>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<3>.NET_005
+ XI1.XI0.XI1<4>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<3>.NET_003
+ XI1.XI0.XI1<4>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_89_4 REG_DATA_4<3> XI1.XI0.XI1<4>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<3>.MM_i_55 XI1.XI0.XI1<4>.XI7<3>.NET_001
+ XI1.XI0.XI1<4>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_61 XI1.XI0.XI1<4>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_66 XI1.XI0.XI1<4>.XI7<3>.NET_003
+ XI1.XI0.XI1<4>.XI7<3>.NET_000 XI1.XI0.XI1<4>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_72 XI1.XI0.XI1<4>.XI7<3>.NET_007
+ XI1.XI0.XI1<4>.XI7<3>.NET_001 XI1.XI0.XI1<4>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<3>.NET_005
+ XI1.XI0.XI1<4>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<3>.NET_003
+ XI1.XI0.XI1<4>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_41_11 REG_DATA_4<2> XI1.XI0.XI1<4>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<2>.MM_i_7 XI1.XI0.XI1<4>.XI7<2>.NET_001
+ XI1.XI0.XI1<4>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_13 XI1.XI0.XI1<4>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_18 XI1.XI0.XI1<4>.XI7<2>.NET_003
+ XI1.XI0.XI1<4>.XI7<2>.NET_001 XI1.XI0.XI1<4>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_24 XI1.XI0.XI1<4>.XI7<2>.NET_004
+ XI1.XI0.XI1<4>.XI7<2>.NET_000 XI1.XI0.XI1<4>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<2>.NET_005
+ XI1.XI0.XI1<4>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<2>.NET_003
+ XI1.XI0.XI1<4>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_89_4 REG_DATA_4<2> XI1.XI0.XI1<4>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<2>.MM_i_55 XI1.XI0.XI1<4>.XI7<2>.NET_001
+ XI1.XI0.XI1<4>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_61 XI1.XI0.XI1<4>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_66 XI1.XI0.XI1<4>.XI7<2>.NET_003
+ XI1.XI0.XI1<4>.XI7<2>.NET_000 XI1.XI0.XI1<4>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_72 XI1.XI0.XI1<4>.XI7<2>.NET_007
+ XI1.XI0.XI1<4>.XI7<2>.NET_001 XI1.XI0.XI1<4>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<2>.NET_005
+ XI1.XI0.XI1<4>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<2>.NET_003
+ XI1.XI0.XI1<4>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_41_11 REG_DATA_4<1> XI1.XI0.XI1<4>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<1>.MM_i_7 XI1.XI0.XI1<4>.XI7<1>.NET_001
+ XI1.XI0.XI1<4>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_13 XI1.XI0.XI1<4>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_18 XI1.XI0.XI1<4>.XI7<1>.NET_003
+ XI1.XI0.XI1<4>.XI7<1>.NET_001 XI1.XI0.XI1<4>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_24 XI1.XI0.XI1<4>.XI7<1>.NET_004
+ XI1.XI0.XI1<4>.XI7<1>.NET_000 XI1.XI0.XI1<4>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<1>.NET_005
+ XI1.XI0.XI1<4>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<1>.NET_003
+ XI1.XI0.XI1<4>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_89_4 REG_DATA_4<1> XI1.XI0.XI1<4>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<1>.MM_i_55 XI1.XI0.XI1<4>.XI7<1>.NET_001
+ XI1.XI0.XI1<4>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_61 XI1.XI0.XI1<4>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_66 XI1.XI0.XI1<4>.XI7<1>.NET_003
+ XI1.XI0.XI1<4>.XI7<1>.NET_000 XI1.XI0.XI1<4>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_72 XI1.XI0.XI1<4>.XI7<1>.NET_007
+ XI1.XI0.XI1<4>.XI7<1>.NET_001 XI1.XI0.XI1<4>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<1>.NET_005
+ XI1.XI0.XI1<4>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<1>.NET_003
+ XI1.XI0.XI1<4>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_41_11 REG_DATA_4<0> XI1.XI0.XI1<4>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<0>.MM_i_7 XI1.XI0.XI1<4>.XI7<0>.NET_001
+ XI1.XI0.XI1<4>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_13 XI1.XI0.XI1<4>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_18 XI1.XI0.XI1<4>.XI7<0>.NET_003
+ XI1.XI0.XI1<4>.XI7<0>.NET_001 XI1.XI0.XI1<4>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_24 XI1.XI0.XI1<4>.XI7<0>.NET_004
+ XI1.XI0.XI1<4>.XI7<0>.NET_000 XI1.XI0.XI1<4>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<0>.NET_005
+ XI1.XI0.XI1<4>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<0>.NET_003
+ XI1.XI0.XI1<4>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_89_4 REG_DATA_4<0> XI1.XI0.XI1<4>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<0>.MM_i_55 XI1.XI0.XI1<4>.XI7<0>.NET_001
+ XI1.XI0.XI1<4>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_61 XI1.XI0.XI1<4>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_66 XI1.XI0.XI1<4>.XI7<0>.NET_003
+ XI1.XI0.XI1<4>.XI7<0>.NET_000 XI1.XI0.XI1<4>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_72 XI1.XI0.XI1<4>.XI7<0>.NET_007
+ XI1.XI0.XI1<4>.XI7<0>.NET_001 XI1.XI0.XI1<4>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<0>.NET_005
+ XI1.XI0.XI1<4>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<0>.NET_003
+ XI1.XI0.XI1<4>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_41_11 REG_DATA_4<7> XI1.XI0.XI1<4>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<7>.MM_i_7 XI1.XI0.XI1<4>.XI7<7>.NET_001
+ XI1.XI0.XI1<4>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_13 XI1.XI0.XI1<4>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_18 XI1.XI0.XI1<4>.XI7<7>.NET_003
+ XI1.XI0.XI1<4>.XI7<7>.NET_001 XI1.XI0.XI1<4>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_24 XI1.XI0.XI1<4>.XI7<7>.NET_004
+ XI1.XI0.XI1<4>.XI7<7>.NET_000 XI1.XI0.XI1<4>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<7>.NET_005
+ XI1.XI0.XI1<4>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<7>.NET_003
+ XI1.XI0.XI1<4>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_89_4 REG_DATA_4<7> XI1.XI0.XI1<4>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<7>.MM_i_55 XI1.XI0.XI1<4>.XI7<7>.NET_001
+ XI1.XI0.XI1<4>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_61 XI1.XI0.XI1<4>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_66 XI1.XI0.XI1<4>.XI7<7>.NET_003
+ XI1.XI0.XI1<4>.XI7<7>.NET_000 XI1.XI0.XI1<4>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_72 XI1.XI0.XI1<4>.XI7<7>.NET_007
+ XI1.XI0.XI1<4>.XI7<7>.NET_001 XI1.XI0.XI1<4>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<7>.NET_005
+ XI1.XI0.XI1<4>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<7>.NET_003
+ XI1.XI0.XI1<4>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_41_11 REG_DATA_4<6> XI1.XI0.XI1<4>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<6>.MM_i_7 XI1.XI0.XI1<4>.XI7<6>.NET_001
+ XI1.XI0.XI1<4>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_13 XI1.XI0.XI1<4>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_18 XI1.XI0.XI1<4>.XI7<6>.NET_003
+ XI1.XI0.XI1<4>.XI7<6>.NET_001 XI1.XI0.XI1<4>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_24 XI1.XI0.XI1<4>.XI7<6>.NET_004
+ XI1.XI0.XI1<4>.XI7<6>.NET_000 XI1.XI0.XI1<4>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<6>.NET_005
+ XI1.XI0.XI1<4>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<6>.NET_003
+ XI1.XI0.XI1<4>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_89_4 REG_DATA_4<6> XI1.XI0.XI1<4>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<6>.MM_i_55 XI1.XI0.XI1<4>.XI7<6>.NET_001
+ XI1.XI0.XI1<4>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_61 XI1.XI0.XI1<4>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_66 XI1.XI0.XI1<4>.XI7<6>.NET_003
+ XI1.XI0.XI1<4>.XI7<6>.NET_000 XI1.XI0.XI1<4>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_72 XI1.XI0.XI1<4>.XI7<6>.NET_007
+ XI1.XI0.XI1<4>.XI7<6>.NET_001 XI1.XI0.XI1<4>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<6>.NET_005
+ XI1.XI0.XI1<4>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<6>.NET_003
+ XI1.XI0.XI1<4>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_41_11 REG_DATA_4<5> XI1.XI0.XI1<4>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<5>.MM_i_7 XI1.XI0.XI1<4>.XI7<5>.NET_001
+ XI1.XI0.XI1<4>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_13 XI1.XI0.XI1<4>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_18 XI1.XI0.XI1<4>.XI7<5>.NET_003
+ XI1.XI0.XI1<4>.XI7<5>.NET_001 XI1.XI0.XI1<4>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_24 XI1.XI0.XI1<4>.XI7<5>.NET_004
+ XI1.XI0.XI1<4>.XI7<5>.NET_000 XI1.XI0.XI1<4>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<5>.NET_005
+ XI1.XI0.XI1<4>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<5>.NET_003
+ XI1.XI0.XI1<4>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_89_4 REG_DATA_4<5> XI1.XI0.XI1<4>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<5>.MM_i_55 XI1.XI0.XI1<4>.XI7<5>.NET_001
+ XI1.XI0.XI1<4>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_61 XI1.XI0.XI1<4>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_66 XI1.XI0.XI1<4>.XI7<5>.NET_003
+ XI1.XI0.XI1<4>.XI7<5>.NET_000 XI1.XI0.XI1<4>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_72 XI1.XI0.XI1<4>.XI7<5>.NET_007
+ XI1.XI0.XI1<4>.XI7<5>.NET_001 XI1.XI0.XI1<4>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<5>.NET_005
+ XI1.XI0.XI1<4>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<5>.NET_003
+ XI1.XI0.XI1<4>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_41_11 REG_DATA_4<4> XI1.XI0.XI1<4>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<4>.MM_i_7 XI1.XI0.XI1<4>.XI7<4>.NET_001
+ XI1.XI0.XI1<4>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_13 XI1.XI0.XI1<4>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_18 XI1.XI0.XI1<4>.XI7<4>.NET_003
+ XI1.XI0.XI1<4>.XI7<4>.NET_001 XI1.XI0.XI1<4>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_24 XI1.XI0.XI1<4>.XI7<4>.NET_004
+ XI1.XI0.XI1<4>.XI7<4>.NET_000 XI1.XI0.XI1<4>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<4>.NET_005
+ XI1.XI0.XI1<4>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<4>.NET_003
+ XI1.XI0.XI1<4>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_89_4 REG_DATA_4<4> XI1.XI0.XI1<4>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<4>.MM_i_55 XI1.XI0.XI1<4>.XI7<4>.NET_001
+ XI1.XI0.XI1<4>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_61 XI1.XI0.XI1<4>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_66 XI1.XI0.XI1<4>.XI7<4>.NET_003
+ XI1.XI0.XI1<4>.XI7<4>.NET_000 XI1.XI0.XI1<4>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_72 XI1.XI0.XI1<4>.XI7<4>.NET_007
+ XI1.XI0.XI1<4>.XI7<4>.NET_001 XI1.XI0.XI1<4>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<4>.NET_005
+ XI1.XI0.XI1<4>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<4>.NET_003
+ XI1.XI0.XI1<4>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_41_11 REG_DATA_4<11> XI1.XI0.XI1<4>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<11>.MM_i_7 XI1.XI0.XI1<4>.XI7<11>.NET_001
+ XI1.XI0.XI1<4>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_13 XI1.XI0.XI1<4>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_18 XI1.XI0.XI1<4>.XI7<11>.NET_003
+ XI1.XI0.XI1<4>.XI7<11>.NET_001 XI1.XI0.XI1<4>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_24 XI1.XI0.XI1<4>.XI7<11>.NET_004
+ XI1.XI0.XI1<4>.XI7<11>.NET_000 XI1.XI0.XI1<4>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<11>.NET_005
+ XI1.XI0.XI1<4>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<11>.NET_003
+ XI1.XI0.XI1<4>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_89_4 REG_DATA_4<11> XI1.XI0.XI1<4>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<11>.MM_i_55 XI1.XI0.XI1<4>.XI7<11>.NET_001
+ XI1.XI0.XI1<4>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_61 XI1.XI0.XI1<4>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_66 XI1.XI0.XI1<4>.XI7<11>.NET_003
+ XI1.XI0.XI1<4>.XI7<11>.NET_000 XI1.XI0.XI1<4>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_72 XI1.XI0.XI1<4>.XI7<11>.NET_007
+ XI1.XI0.XI1<4>.XI7<11>.NET_001 XI1.XI0.XI1<4>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<11>.NET_005
+ XI1.XI0.XI1<4>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<11>.NET_003
+ XI1.XI0.XI1<4>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_41_11 REG_DATA_4<10> XI1.XI0.XI1<4>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<10>.MM_i_7 XI1.XI0.XI1<4>.XI7<10>.NET_001
+ XI1.XI0.XI1<4>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_13 XI1.XI0.XI1<4>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_18 XI1.XI0.XI1<4>.XI7<10>.NET_003
+ XI1.XI0.XI1<4>.XI7<10>.NET_001 XI1.XI0.XI1<4>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_24 XI1.XI0.XI1<4>.XI7<10>.NET_004
+ XI1.XI0.XI1<4>.XI7<10>.NET_000 XI1.XI0.XI1<4>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<10>.NET_005
+ XI1.XI0.XI1<4>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<10>.NET_003
+ XI1.XI0.XI1<4>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_89_4 REG_DATA_4<10> XI1.XI0.XI1<4>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<10>.MM_i_55 XI1.XI0.XI1<4>.XI7<10>.NET_001
+ XI1.XI0.XI1<4>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_61 XI1.XI0.XI1<4>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_66 XI1.XI0.XI1<4>.XI7<10>.NET_003
+ XI1.XI0.XI1<4>.XI7<10>.NET_000 XI1.XI0.XI1<4>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_72 XI1.XI0.XI1<4>.XI7<10>.NET_007
+ XI1.XI0.XI1<4>.XI7<10>.NET_001 XI1.XI0.XI1<4>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<10>.NET_005
+ XI1.XI0.XI1<4>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<10>.NET_003
+ XI1.XI0.XI1<4>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_41_11 REG_DATA_4<9> XI1.XI0.XI1<4>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<9>.MM_i_7 XI1.XI0.XI1<4>.XI7<9>.NET_001
+ XI1.XI0.XI1<4>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_13 XI1.XI0.XI1<4>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_18 XI1.XI0.XI1<4>.XI7<9>.NET_003
+ XI1.XI0.XI1<4>.XI7<9>.NET_001 XI1.XI0.XI1<4>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_24 XI1.XI0.XI1<4>.XI7<9>.NET_004
+ XI1.XI0.XI1<4>.XI7<9>.NET_000 XI1.XI0.XI1<4>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<9>.NET_005
+ XI1.XI0.XI1<4>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<9>.NET_003
+ XI1.XI0.XI1<4>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_89_4 REG_DATA_4<9> XI1.XI0.XI1<4>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<9>.MM_i_55 XI1.XI0.XI1<4>.XI7<9>.NET_001
+ XI1.XI0.XI1<4>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_61 XI1.XI0.XI1<4>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_66 XI1.XI0.XI1<4>.XI7<9>.NET_003
+ XI1.XI0.XI1<4>.XI7<9>.NET_000 XI1.XI0.XI1<4>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_72 XI1.XI0.XI1<4>.XI7<9>.NET_007
+ XI1.XI0.XI1<4>.XI7<9>.NET_001 XI1.XI0.XI1<4>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<9>.NET_005
+ XI1.XI0.XI1<4>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<9>.NET_003
+ XI1.XI0.XI1<4>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_41_11 REG_DATA_4<8> XI1.XI0.XI1<4>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<8>.MM_i_7 XI1.XI0.XI1<4>.XI7<8>.NET_001
+ XI1.XI0.XI1<4>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_13 XI1.XI0.XI1<4>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_18 XI1.XI0.XI1<4>.XI7<8>.NET_003
+ XI1.XI0.XI1<4>.XI7<8>.NET_001 XI1.XI0.XI1<4>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_24 XI1.XI0.XI1<4>.XI7<8>.NET_004
+ XI1.XI0.XI1<4>.XI7<8>.NET_000 XI1.XI0.XI1<4>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<8>.NET_005
+ XI1.XI0.XI1<4>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<8>.NET_003
+ XI1.XI0.XI1<4>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_89_4 REG_DATA_4<8> XI1.XI0.XI1<4>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<8>.MM_i_55 XI1.XI0.XI1<4>.XI7<8>.NET_001
+ XI1.XI0.XI1<4>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_61 XI1.XI0.XI1<4>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_66 XI1.XI0.XI1<4>.XI7<8>.NET_003
+ XI1.XI0.XI1<4>.XI7<8>.NET_000 XI1.XI0.XI1<4>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_72 XI1.XI0.XI1<4>.XI7<8>.NET_007
+ XI1.XI0.XI1<4>.XI7<8>.NET_001 XI1.XI0.XI1<4>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<8>.NET_005
+ XI1.XI0.XI1<4>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<8>.NET_003
+ XI1.XI0.XI1<4>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_41_11 REG_DATA_4<15> XI1.XI0.XI1<4>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<15>.MM_i_7 XI1.XI0.XI1<4>.XI7<15>.NET_001
+ XI1.XI0.XI1<4>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_13 XI1.XI0.XI1<4>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_18 XI1.XI0.XI1<4>.XI7<15>.NET_003
+ XI1.XI0.XI1<4>.XI7<15>.NET_001 XI1.XI0.XI1<4>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_24 XI1.XI0.XI1<4>.XI7<15>.NET_004
+ XI1.XI0.XI1<4>.XI7<15>.NET_000 XI1.XI0.XI1<4>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<15>.NET_005
+ XI1.XI0.XI1<4>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<15>.NET_003
+ XI1.XI0.XI1<4>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_89_4 REG_DATA_4<15> XI1.XI0.XI1<4>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<15>.MM_i_55 XI1.XI0.XI1<4>.XI7<15>.NET_001
+ XI1.XI0.XI1<4>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_61 XI1.XI0.XI1<4>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_66 XI1.XI0.XI1<4>.XI7<15>.NET_003
+ XI1.XI0.XI1<4>.XI7<15>.NET_000 XI1.XI0.XI1<4>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_72 XI1.XI0.XI1<4>.XI7<15>.NET_007
+ XI1.XI0.XI1<4>.XI7<15>.NET_001 XI1.XI0.XI1<4>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<15>.NET_005
+ XI1.XI0.XI1<4>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<15>.NET_003
+ XI1.XI0.XI1<4>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_41_11 REG_DATA_4<14> XI1.XI0.XI1<4>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<14>.MM_i_7 XI1.XI0.XI1<4>.XI7<14>.NET_001
+ XI1.XI0.XI1<4>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_13 XI1.XI0.XI1<4>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_18 XI1.XI0.XI1<4>.XI7<14>.NET_003
+ XI1.XI0.XI1<4>.XI7<14>.NET_001 XI1.XI0.XI1<4>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_24 XI1.XI0.XI1<4>.XI7<14>.NET_004
+ XI1.XI0.XI1<4>.XI7<14>.NET_000 XI1.XI0.XI1<4>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<14>.NET_005
+ XI1.XI0.XI1<4>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<14>.NET_003
+ XI1.XI0.XI1<4>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_89_4 REG_DATA_4<14> XI1.XI0.XI1<4>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<14>.MM_i_55 XI1.XI0.XI1<4>.XI7<14>.NET_001
+ XI1.XI0.XI1<4>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_61 XI1.XI0.XI1<4>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_66 XI1.XI0.XI1<4>.XI7<14>.NET_003
+ XI1.XI0.XI1<4>.XI7<14>.NET_000 XI1.XI0.XI1<4>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_72 XI1.XI0.XI1<4>.XI7<14>.NET_007
+ XI1.XI0.XI1<4>.XI7<14>.NET_001 XI1.XI0.XI1<4>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<14>.NET_005
+ XI1.XI0.XI1<4>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<14>.NET_003
+ XI1.XI0.XI1<4>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_41_11 REG_DATA_4<13> XI1.XI0.XI1<4>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<13>.MM_i_7 XI1.XI0.XI1<4>.XI7<13>.NET_001
+ XI1.XI0.XI1<4>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_13 XI1.XI0.XI1<4>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_18 XI1.XI0.XI1<4>.XI7<13>.NET_003
+ XI1.XI0.XI1<4>.XI7<13>.NET_001 XI1.XI0.XI1<4>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_24 XI1.XI0.XI1<4>.XI7<13>.NET_004
+ XI1.XI0.XI1<4>.XI7<13>.NET_000 XI1.XI0.XI1<4>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<13>.NET_005
+ XI1.XI0.XI1<4>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<13>.NET_003
+ XI1.XI0.XI1<4>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_89_4 REG_DATA_4<13> XI1.XI0.XI1<4>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<13>.MM_i_55 XI1.XI0.XI1<4>.XI7<13>.NET_001
+ XI1.XI0.XI1<4>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_61 XI1.XI0.XI1<4>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_66 XI1.XI0.XI1<4>.XI7<13>.NET_003
+ XI1.XI0.XI1<4>.XI7<13>.NET_000 XI1.XI0.XI1<4>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_72 XI1.XI0.XI1<4>.XI7<13>.NET_007
+ XI1.XI0.XI1<4>.XI7<13>.NET_001 XI1.XI0.XI1<4>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<13>.NET_005
+ XI1.XI0.XI1<4>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<13>.NET_003
+ XI1.XI0.XI1<4>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_41_11 REG_DATA_4<12> XI1.XI0.XI1<4>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<4>.XI7<12>.MM_i_7 XI1.XI0.XI1<4>.XI7<12>.NET_001
+ XI1.XI0.XI1<4>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_13 XI1.XI0.XI1<4>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_18 XI1.XI0.XI1<4>.XI7<12>.NET_003
+ XI1.XI0.XI1<4>.XI7<12>.NET_001 XI1.XI0.XI1<4>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_24 XI1.XI0.XI1<4>.XI7<12>.NET_004
+ XI1.XI0.XI1<4>.XI7<12>.NET_000 XI1.XI0.XI1<4>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<4>.XI7<12>.NET_005
+ XI1.XI0.XI1<4>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<4>.XI7<12>.NET_003
+ XI1.XI0.XI1<4>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<4>
+ XI1.XI0.XI1<4>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_89_4 REG_DATA_4<12> XI1.XI0.XI1<4>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<4>.XI7<12>.MM_i_55 XI1.XI0.XI1<4>.XI7<12>.NET_001
+ XI1.XI0.XI1<4>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_61 XI1.XI0.XI1<4>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_66 XI1.XI0.XI1<4>.XI7<12>.NET_003
+ XI1.XI0.XI1<4>.XI7<12>.NET_000 XI1.XI0.XI1<4>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_72 XI1.XI0.XI1<4>.XI7<12>.NET_007
+ XI1.XI0.XI1<4>.XI7<12>.NET_001 XI1.XI0.XI1<4>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<4>.XI7<12>.NET_005
+ XI1.XI0.XI1<4>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<4>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<4>.XI7<12>.NET_003
+ XI1.XI0.XI1<4>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_41_11 REG_DATA_3<3> XI1.XI0.XI1<3>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<3>.MM_i_7 XI1.XI0.XI1<3>.XI7<3>.NET_001
+ XI1.XI0.XI1<3>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_13 XI1.XI0.XI1<3>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_18 XI1.XI0.XI1<3>.XI7<3>.NET_003
+ XI1.XI0.XI1<3>.XI7<3>.NET_001 XI1.XI0.XI1<3>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_24 XI1.XI0.XI1<3>.XI7<3>.NET_004
+ XI1.XI0.XI1<3>.XI7<3>.NET_000 XI1.XI0.XI1<3>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<3>.NET_005
+ XI1.XI0.XI1<3>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<3>.NET_003
+ XI1.XI0.XI1<3>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_89_4 REG_DATA_3<3> XI1.XI0.XI1<3>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<3>.MM_i_55 XI1.XI0.XI1<3>.XI7<3>.NET_001
+ XI1.XI0.XI1<3>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_61 XI1.XI0.XI1<3>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_66 XI1.XI0.XI1<3>.XI7<3>.NET_003
+ XI1.XI0.XI1<3>.XI7<3>.NET_000 XI1.XI0.XI1<3>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_72 XI1.XI0.XI1<3>.XI7<3>.NET_007
+ XI1.XI0.XI1<3>.XI7<3>.NET_001 XI1.XI0.XI1<3>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<3>.NET_005
+ XI1.XI0.XI1<3>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<3>.NET_003
+ XI1.XI0.XI1<3>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_41_11 REG_DATA_3<2> XI1.XI0.XI1<3>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<2>.MM_i_7 XI1.XI0.XI1<3>.XI7<2>.NET_001
+ XI1.XI0.XI1<3>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_13 XI1.XI0.XI1<3>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_18 XI1.XI0.XI1<3>.XI7<2>.NET_003
+ XI1.XI0.XI1<3>.XI7<2>.NET_001 XI1.XI0.XI1<3>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_24 XI1.XI0.XI1<3>.XI7<2>.NET_004
+ XI1.XI0.XI1<3>.XI7<2>.NET_000 XI1.XI0.XI1<3>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<2>.NET_005
+ XI1.XI0.XI1<3>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<2>.NET_003
+ XI1.XI0.XI1<3>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_89_4 REG_DATA_3<2> XI1.XI0.XI1<3>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<2>.MM_i_55 XI1.XI0.XI1<3>.XI7<2>.NET_001
+ XI1.XI0.XI1<3>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_61 XI1.XI0.XI1<3>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_66 XI1.XI0.XI1<3>.XI7<2>.NET_003
+ XI1.XI0.XI1<3>.XI7<2>.NET_000 XI1.XI0.XI1<3>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_72 XI1.XI0.XI1<3>.XI7<2>.NET_007
+ XI1.XI0.XI1<3>.XI7<2>.NET_001 XI1.XI0.XI1<3>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<2>.NET_005
+ XI1.XI0.XI1<3>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<2>.NET_003
+ XI1.XI0.XI1<3>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_41_11 REG_DATA_3<1> XI1.XI0.XI1<3>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<1>.MM_i_7 XI1.XI0.XI1<3>.XI7<1>.NET_001
+ XI1.XI0.XI1<3>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_13 XI1.XI0.XI1<3>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_18 XI1.XI0.XI1<3>.XI7<1>.NET_003
+ XI1.XI0.XI1<3>.XI7<1>.NET_001 XI1.XI0.XI1<3>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_24 XI1.XI0.XI1<3>.XI7<1>.NET_004
+ XI1.XI0.XI1<3>.XI7<1>.NET_000 XI1.XI0.XI1<3>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<1>.NET_005
+ XI1.XI0.XI1<3>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<1>.NET_003
+ XI1.XI0.XI1<3>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_89_4 REG_DATA_3<1> XI1.XI0.XI1<3>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<1>.MM_i_55 XI1.XI0.XI1<3>.XI7<1>.NET_001
+ XI1.XI0.XI1<3>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_61 XI1.XI0.XI1<3>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_66 XI1.XI0.XI1<3>.XI7<1>.NET_003
+ XI1.XI0.XI1<3>.XI7<1>.NET_000 XI1.XI0.XI1<3>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_72 XI1.XI0.XI1<3>.XI7<1>.NET_007
+ XI1.XI0.XI1<3>.XI7<1>.NET_001 XI1.XI0.XI1<3>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<1>.NET_005
+ XI1.XI0.XI1<3>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<1>.NET_003
+ XI1.XI0.XI1<3>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_41_11 REG_DATA_3<0> XI1.XI0.XI1<3>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<0>.MM_i_7 XI1.XI0.XI1<3>.XI7<0>.NET_001
+ XI1.XI0.XI1<3>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_13 XI1.XI0.XI1<3>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_18 XI1.XI0.XI1<3>.XI7<0>.NET_003
+ XI1.XI0.XI1<3>.XI7<0>.NET_001 XI1.XI0.XI1<3>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_24 XI1.XI0.XI1<3>.XI7<0>.NET_004
+ XI1.XI0.XI1<3>.XI7<0>.NET_000 XI1.XI0.XI1<3>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<0>.NET_005
+ XI1.XI0.XI1<3>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<0>.NET_003
+ XI1.XI0.XI1<3>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_89_4 REG_DATA_3<0> XI1.XI0.XI1<3>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<0>.MM_i_55 XI1.XI0.XI1<3>.XI7<0>.NET_001
+ XI1.XI0.XI1<3>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_61 XI1.XI0.XI1<3>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_66 XI1.XI0.XI1<3>.XI7<0>.NET_003
+ XI1.XI0.XI1<3>.XI7<0>.NET_000 XI1.XI0.XI1<3>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_72 XI1.XI0.XI1<3>.XI7<0>.NET_007
+ XI1.XI0.XI1<3>.XI7<0>.NET_001 XI1.XI0.XI1<3>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<0>.NET_005
+ XI1.XI0.XI1<3>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<0>.NET_003
+ XI1.XI0.XI1<3>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_41_11 REG_DATA_3<7> XI1.XI0.XI1<3>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<7>.MM_i_7 XI1.XI0.XI1<3>.XI7<7>.NET_001
+ XI1.XI0.XI1<3>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_13 XI1.XI0.XI1<3>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_18 XI1.XI0.XI1<3>.XI7<7>.NET_003
+ XI1.XI0.XI1<3>.XI7<7>.NET_001 XI1.XI0.XI1<3>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_24 XI1.XI0.XI1<3>.XI7<7>.NET_004
+ XI1.XI0.XI1<3>.XI7<7>.NET_000 XI1.XI0.XI1<3>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<7>.NET_005
+ XI1.XI0.XI1<3>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<7>.NET_003
+ XI1.XI0.XI1<3>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_89_4 REG_DATA_3<7> XI1.XI0.XI1<3>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<7>.MM_i_55 XI1.XI0.XI1<3>.XI7<7>.NET_001
+ XI1.XI0.XI1<3>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_61 XI1.XI0.XI1<3>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_66 XI1.XI0.XI1<3>.XI7<7>.NET_003
+ XI1.XI0.XI1<3>.XI7<7>.NET_000 XI1.XI0.XI1<3>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_72 XI1.XI0.XI1<3>.XI7<7>.NET_007
+ XI1.XI0.XI1<3>.XI7<7>.NET_001 XI1.XI0.XI1<3>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<7>.NET_005
+ XI1.XI0.XI1<3>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<7>.NET_003
+ XI1.XI0.XI1<3>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_41_11 REG_DATA_3<6> XI1.XI0.XI1<3>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<6>.MM_i_7 XI1.XI0.XI1<3>.XI7<6>.NET_001
+ XI1.XI0.XI1<3>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_13 XI1.XI0.XI1<3>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_18 XI1.XI0.XI1<3>.XI7<6>.NET_003
+ XI1.XI0.XI1<3>.XI7<6>.NET_001 XI1.XI0.XI1<3>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_24 XI1.XI0.XI1<3>.XI7<6>.NET_004
+ XI1.XI0.XI1<3>.XI7<6>.NET_000 XI1.XI0.XI1<3>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<6>.NET_005
+ XI1.XI0.XI1<3>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<6>.NET_003
+ XI1.XI0.XI1<3>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_89_4 REG_DATA_3<6> XI1.XI0.XI1<3>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<6>.MM_i_55 XI1.XI0.XI1<3>.XI7<6>.NET_001
+ XI1.XI0.XI1<3>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_61 XI1.XI0.XI1<3>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_66 XI1.XI0.XI1<3>.XI7<6>.NET_003
+ XI1.XI0.XI1<3>.XI7<6>.NET_000 XI1.XI0.XI1<3>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_72 XI1.XI0.XI1<3>.XI7<6>.NET_007
+ XI1.XI0.XI1<3>.XI7<6>.NET_001 XI1.XI0.XI1<3>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<6>.NET_005
+ XI1.XI0.XI1<3>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<6>.NET_003
+ XI1.XI0.XI1<3>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_41_11 REG_DATA_3<5> XI1.XI0.XI1<3>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<5>.MM_i_7 XI1.XI0.XI1<3>.XI7<5>.NET_001
+ XI1.XI0.XI1<3>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_13 XI1.XI0.XI1<3>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_18 XI1.XI0.XI1<3>.XI7<5>.NET_003
+ XI1.XI0.XI1<3>.XI7<5>.NET_001 XI1.XI0.XI1<3>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_24 XI1.XI0.XI1<3>.XI7<5>.NET_004
+ XI1.XI0.XI1<3>.XI7<5>.NET_000 XI1.XI0.XI1<3>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<5>.NET_005
+ XI1.XI0.XI1<3>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<5>.NET_003
+ XI1.XI0.XI1<3>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_89_4 REG_DATA_3<5> XI1.XI0.XI1<3>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<5>.MM_i_55 XI1.XI0.XI1<3>.XI7<5>.NET_001
+ XI1.XI0.XI1<3>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_61 XI1.XI0.XI1<3>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_66 XI1.XI0.XI1<3>.XI7<5>.NET_003
+ XI1.XI0.XI1<3>.XI7<5>.NET_000 XI1.XI0.XI1<3>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_72 XI1.XI0.XI1<3>.XI7<5>.NET_007
+ XI1.XI0.XI1<3>.XI7<5>.NET_001 XI1.XI0.XI1<3>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<5>.NET_005
+ XI1.XI0.XI1<3>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<5>.NET_003
+ XI1.XI0.XI1<3>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_41_11 REG_DATA_3<4> XI1.XI0.XI1<3>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<4>.MM_i_7 XI1.XI0.XI1<3>.XI7<4>.NET_001
+ XI1.XI0.XI1<3>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_13 XI1.XI0.XI1<3>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_18 XI1.XI0.XI1<3>.XI7<4>.NET_003
+ XI1.XI0.XI1<3>.XI7<4>.NET_001 XI1.XI0.XI1<3>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_24 XI1.XI0.XI1<3>.XI7<4>.NET_004
+ XI1.XI0.XI1<3>.XI7<4>.NET_000 XI1.XI0.XI1<3>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<4>.NET_005
+ XI1.XI0.XI1<3>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<4>.NET_003
+ XI1.XI0.XI1<3>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_89_4 REG_DATA_3<4> XI1.XI0.XI1<3>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<4>.MM_i_55 XI1.XI0.XI1<3>.XI7<4>.NET_001
+ XI1.XI0.XI1<3>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_61 XI1.XI0.XI1<3>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_66 XI1.XI0.XI1<3>.XI7<4>.NET_003
+ XI1.XI0.XI1<3>.XI7<4>.NET_000 XI1.XI0.XI1<3>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_72 XI1.XI0.XI1<3>.XI7<4>.NET_007
+ XI1.XI0.XI1<3>.XI7<4>.NET_001 XI1.XI0.XI1<3>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<4>.NET_005
+ XI1.XI0.XI1<3>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<4>.NET_003
+ XI1.XI0.XI1<3>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_41_11 REG_DATA_3<11> XI1.XI0.XI1<3>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<11>.MM_i_7 XI1.XI0.XI1<3>.XI7<11>.NET_001
+ XI1.XI0.XI1<3>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_13 XI1.XI0.XI1<3>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_18 XI1.XI0.XI1<3>.XI7<11>.NET_003
+ XI1.XI0.XI1<3>.XI7<11>.NET_001 XI1.XI0.XI1<3>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_24 XI1.XI0.XI1<3>.XI7<11>.NET_004
+ XI1.XI0.XI1<3>.XI7<11>.NET_000 XI1.XI0.XI1<3>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<11>.NET_005
+ XI1.XI0.XI1<3>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<11>.NET_003
+ XI1.XI0.XI1<3>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_89_4 REG_DATA_3<11> XI1.XI0.XI1<3>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<11>.MM_i_55 XI1.XI0.XI1<3>.XI7<11>.NET_001
+ XI1.XI0.XI1<3>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_61 XI1.XI0.XI1<3>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_66 XI1.XI0.XI1<3>.XI7<11>.NET_003
+ XI1.XI0.XI1<3>.XI7<11>.NET_000 XI1.XI0.XI1<3>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_72 XI1.XI0.XI1<3>.XI7<11>.NET_007
+ XI1.XI0.XI1<3>.XI7<11>.NET_001 XI1.XI0.XI1<3>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<11>.NET_005
+ XI1.XI0.XI1<3>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<11>.NET_003
+ XI1.XI0.XI1<3>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_41_11 REG_DATA_3<10> XI1.XI0.XI1<3>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<10>.MM_i_7 XI1.XI0.XI1<3>.XI7<10>.NET_001
+ XI1.XI0.XI1<3>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_13 XI1.XI0.XI1<3>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_18 XI1.XI0.XI1<3>.XI7<10>.NET_003
+ XI1.XI0.XI1<3>.XI7<10>.NET_001 XI1.XI0.XI1<3>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_24 XI1.XI0.XI1<3>.XI7<10>.NET_004
+ XI1.XI0.XI1<3>.XI7<10>.NET_000 XI1.XI0.XI1<3>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<10>.NET_005
+ XI1.XI0.XI1<3>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<10>.NET_003
+ XI1.XI0.XI1<3>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_89_4 REG_DATA_3<10> XI1.XI0.XI1<3>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<10>.MM_i_55 XI1.XI0.XI1<3>.XI7<10>.NET_001
+ XI1.XI0.XI1<3>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_61 XI1.XI0.XI1<3>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_66 XI1.XI0.XI1<3>.XI7<10>.NET_003
+ XI1.XI0.XI1<3>.XI7<10>.NET_000 XI1.XI0.XI1<3>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_72 XI1.XI0.XI1<3>.XI7<10>.NET_007
+ XI1.XI0.XI1<3>.XI7<10>.NET_001 XI1.XI0.XI1<3>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<10>.NET_005
+ XI1.XI0.XI1<3>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<10>.NET_003
+ XI1.XI0.XI1<3>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_41_11 REG_DATA_3<9> XI1.XI0.XI1<3>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<9>.MM_i_7 XI1.XI0.XI1<3>.XI7<9>.NET_001
+ XI1.XI0.XI1<3>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_13 XI1.XI0.XI1<3>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_18 XI1.XI0.XI1<3>.XI7<9>.NET_003
+ XI1.XI0.XI1<3>.XI7<9>.NET_001 XI1.XI0.XI1<3>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_24 XI1.XI0.XI1<3>.XI7<9>.NET_004
+ XI1.XI0.XI1<3>.XI7<9>.NET_000 XI1.XI0.XI1<3>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<9>.NET_005
+ XI1.XI0.XI1<3>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<9>.NET_003
+ XI1.XI0.XI1<3>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_89_4 REG_DATA_3<9> XI1.XI0.XI1<3>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<9>.MM_i_55 XI1.XI0.XI1<3>.XI7<9>.NET_001
+ XI1.XI0.XI1<3>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_61 XI1.XI0.XI1<3>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_66 XI1.XI0.XI1<3>.XI7<9>.NET_003
+ XI1.XI0.XI1<3>.XI7<9>.NET_000 XI1.XI0.XI1<3>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_72 XI1.XI0.XI1<3>.XI7<9>.NET_007
+ XI1.XI0.XI1<3>.XI7<9>.NET_001 XI1.XI0.XI1<3>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<9>.NET_005
+ XI1.XI0.XI1<3>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<9>.NET_003
+ XI1.XI0.XI1<3>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_41_11 REG_DATA_3<8> XI1.XI0.XI1<3>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<8>.MM_i_7 XI1.XI0.XI1<3>.XI7<8>.NET_001
+ XI1.XI0.XI1<3>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_13 XI1.XI0.XI1<3>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_18 XI1.XI0.XI1<3>.XI7<8>.NET_003
+ XI1.XI0.XI1<3>.XI7<8>.NET_001 XI1.XI0.XI1<3>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_24 XI1.XI0.XI1<3>.XI7<8>.NET_004
+ XI1.XI0.XI1<3>.XI7<8>.NET_000 XI1.XI0.XI1<3>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<8>.NET_005
+ XI1.XI0.XI1<3>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<8>.NET_003
+ XI1.XI0.XI1<3>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_89_4 REG_DATA_3<8> XI1.XI0.XI1<3>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<8>.MM_i_55 XI1.XI0.XI1<3>.XI7<8>.NET_001
+ XI1.XI0.XI1<3>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_61 XI1.XI0.XI1<3>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_66 XI1.XI0.XI1<3>.XI7<8>.NET_003
+ XI1.XI0.XI1<3>.XI7<8>.NET_000 XI1.XI0.XI1<3>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_72 XI1.XI0.XI1<3>.XI7<8>.NET_007
+ XI1.XI0.XI1<3>.XI7<8>.NET_001 XI1.XI0.XI1<3>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<8>.NET_005
+ XI1.XI0.XI1<3>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<8>.NET_003
+ XI1.XI0.XI1<3>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_41_11 REG_DATA_3<15> XI1.XI0.XI1<3>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<15>.MM_i_7 XI1.XI0.XI1<3>.XI7<15>.NET_001
+ XI1.XI0.XI1<3>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_13 XI1.XI0.XI1<3>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_18 XI1.XI0.XI1<3>.XI7<15>.NET_003
+ XI1.XI0.XI1<3>.XI7<15>.NET_001 XI1.XI0.XI1<3>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_24 XI1.XI0.XI1<3>.XI7<15>.NET_004
+ XI1.XI0.XI1<3>.XI7<15>.NET_000 XI1.XI0.XI1<3>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<15>.NET_005
+ XI1.XI0.XI1<3>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<15>.NET_003
+ XI1.XI0.XI1<3>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_89_4 REG_DATA_3<15> XI1.XI0.XI1<3>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<15>.MM_i_55 XI1.XI0.XI1<3>.XI7<15>.NET_001
+ XI1.XI0.XI1<3>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_61 XI1.XI0.XI1<3>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_66 XI1.XI0.XI1<3>.XI7<15>.NET_003
+ XI1.XI0.XI1<3>.XI7<15>.NET_000 XI1.XI0.XI1<3>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_72 XI1.XI0.XI1<3>.XI7<15>.NET_007
+ XI1.XI0.XI1<3>.XI7<15>.NET_001 XI1.XI0.XI1<3>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<15>.NET_005
+ XI1.XI0.XI1<3>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<15>.NET_003
+ XI1.XI0.XI1<3>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_41_11 REG_DATA_3<14> XI1.XI0.XI1<3>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<14>.MM_i_7 XI1.XI0.XI1<3>.XI7<14>.NET_001
+ XI1.XI0.XI1<3>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_13 XI1.XI0.XI1<3>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_18 XI1.XI0.XI1<3>.XI7<14>.NET_003
+ XI1.XI0.XI1<3>.XI7<14>.NET_001 XI1.XI0.XI1<3>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_24 XI1.XI0.XI1<3>.XI7<14>.NET_004
+ XI1.XI0.XI1<3>.XI7<14>.NET_000 XI1.XI0.XI1<3>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<14>.NET_005
+ XI1.XI0.XI1<3>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<14>.NET_003
+ XI1.XI0.XI1<3>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_89_4 REG_DATA_3<14> XI1.XI0.XI1<3>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<14>.MM_i_55 XI1.XI0.XI1<3>.XI7<14>.NET_001
+ XI1.XI0.XI1<3>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_61 XI1.XI0.XI1<3>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_66 XI1.XI0.XI1<3>.XI7<14>.NET_003
+ XI1.XI0.XI1<3>.XI7<14>.NET_000 XI1.XI0.XI1<3>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_72 XI1.XI0.XI1<3>.XI7<14>.NET_007
+ XI1.XI0.XI1<3>.XI7<14>.NET_001 XI1.XI0.XI1<3>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<14>.NET_005
+ XI1.XI0.XI1<3>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<14>.NET_003
+ XI1.XI0.XI1<3>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_41_11 REG_DATA_3<13> XI1.XI0.XI1<3>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<13>.MM_i_7 XI1.XI0.XI1<3>.XI7<13>.NET_001
+ XI1.XI0.XI1<3>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_13 XI1.XI0.XI1<3>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_18 XI1.XI0.XI1<3>.XI7<13>.NET_003
+ XI1.XI0.XI1<3>.XI7<13>.NET_001 XI1.XI0.XI1<3>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_24 XI1.XI0.XI1<3>.XI7<13>.NET_004
+ XI1.XI0.XI1<3>.XI7<13>.NET_000 XI1.XI0.XI1<3>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<13>.NET_005
+ XI1.XI0.XI1<3>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<13>.NET_003
+ XI1.XI0.XI1<3>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_89_4 REG_DATA_3<13> XI1.XI0.XI1<3>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<13>.MM_i_55 XI1.XI0.XI1<3>.XI7<13>.NET_001
+ XI1.XI0.XI1<3>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_61 XI1.XI0.XI1<3>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_66 XI1.XI0.XI1<3>.XI7<13>.NET_003
+ XI1.XI0.XI1<3>.XI7<13>.NET_000 XI1.XI0.XI1<3>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_72 XI1.XI0.XI1<3>.XI7<13>.NET_007
+ XI1.XI0.XI1<3>.XI7<13>.NET_001 XI1.XI0.XI1<3>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<13>.NET_005
+ XI1.XI0.XI1<3>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<13>.NET_003
+ XI1.XI0.XI1<3>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_41_11 REG_DATA_3<12> XI1.XI0.XI1<3>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<3>.XI7<12>.MM_i_7 XI1.XI0.XI1<3>.XI7<12>.NET_001
+ XI1.XI0.XI1<3>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_13 XI1.XI0.XI1<3>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_18 XI1.XI0.XI1<3>.XI7<12>.NET_003
+ XI1.XI0.XI1<3>.XI7<12>.NET_001 XI1.XI0.XI1<3>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_24 XI1.XI0.XI1<3>.XI7<12>.NET_004
+ XI1.XI0.XI1<3>.XI7<12>.NET_000 XI1.XI0.XI1<3>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<3>.XI7<12>.NET_005
+ XI1.XI0.XI1<3>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<3>.XI7<12>.NET_003
+ XI1.XI0.XI1<3>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<3>
+ XI1.XI0.XI1<3>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_89_4 REG_DATA_3<12> XI1.XI0.XI1<3>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<3>.XI7<12>.MM_i_55 XI1.XI0.XI1<3>.XI7<12>.NET_001
+ XI1.XI0.XI1<3>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_61 XI1.XI0.XI1<3>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_66 XI1.XI0.XI1<3>.XI7<12>.NET_003
+ XI1.XI0.XI1<3>.XI7<12>.NET_000 XI1.XI0.XI1<3>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_72 XI1.XI0.XI1<3>.XI7<12>.NET_007
+ XI1.XI0.XI1<3>.XI7<12>.NET_001 XI1.XI0.XI1<3>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<3>.XI7<12>.NET_005
+ XI1.XI0.XI1<3>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<3>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<3>.XI7<12>.NET_003
+ XI1.XI0.XI1<3>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_41_11 REG_DATA_2<3> XI1.XI0.XI1<2>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<3>.MM_i_7 XI1.XI0.XI1<2>.XI7<3>.NET_001
+ XI1.XI0.XI1<2>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_13 XI1.XI0.XI1<2>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_18 XI1.XI0.XI1<2>.XI7<3>.NET_003
+ XI1.XI0.XI1<2>.XI7<3>.NET_001 XI1.XI0.XI1<2>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_24 XI1.XI0.XI1<2>.XI7<3>.NET_004
+ XI1.XI0.XI1<2>.XI7<3>.NET_000 XI1.XI0.XI1<2>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<3>.NET_005
+ XI1.XI0.XI1<2>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<3>.NET_003
+ XI1.XI0.XI1<2>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_89_4 REG_DATA_2<3> XI1.XI0.XI1<2>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<3>.MM_i_55 XI1.XI0.XI1<2>.XI7<3>.NET_001
+ XI1.XI0.XI1<2>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_61 XI1.XI0.XI1<2>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_66 XI1.XI0.XI1<2>.XI7<3>.NET_003
+ XI1.XI0.XI1<2>.XI7<3>.NET_000 XI1.XI0.XI1<2>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_72 XI1.XI0.XI1<2>.XI7<3>.NET_007
+ XI1.XI0.XI1<2>.XI7<3>.NET_001 XI1.XI0.XI1<2>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<3>.NET_005
+ XI1.XI0.XI1<2>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<3>.NET_003
+ XI1.XI0.XI1<2>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_41_11 REG_DATA_2<2> XI1.XI0.XI1<2>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<2>.MM_i_7 XI1.XI0.XI1<2>.XI7<2>.NET_001
+ XI1.XI0.XI1<2>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_13 XI1.XI0.XI1<2>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_18 XI1.XI0.XI1<2>.XI7<2>.NET_003
+ XI1.XI0.XI1<2>.XI7<2>.NET_001 XI1.XI0.XI1<2>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_24 XI1.XI0.XI1<2>.XI7<2>.NET_004
+ XI1.XI0.XI1<2>.XI7<2>.NET_000 XI1.XI0.XI1<2>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<2>.NET_005
+ XI1.XI0.XI1<2>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<2>.NET_003
+ XI1.XI0.XI1<2>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_89_4 REG_DATA_2<2> XI1.XI0.XI1<2>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<2>.MM_i_55 XI1.XI0.XI1<2>.XI7<2>.NET_001
+ XI1.XI0.XI1<2>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_61 XI1.XI0.XI1<2>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_66 XI1.XI0.XI1<2>.XI7<2>.NET_003
+ XI1.XI0.XI1<2>.XI7<2>.NET_000 XI1.XI0.XI1<2>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_72 XI1.XI0.XI1<2>.XI7<2>.NET_007
+ XI1.XI0.XI1<2>.XI7<2>.NET_001 XI1.XI0.XI1<2>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<2>.NET_005
+ XI1.XI0.XI1<2>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<2>.NET_003
+ XI1.XI0.XI1<2>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_41_11 REG_DATA_2<1> XI1.XI0.XI1<2>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<1>.MM_i_7 XI1.XI0.XI1<2>.XI7<1>.NET_001
+ XI1.XI0.XI1<2>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_13 XI1.XI0.XI1<2>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_18 XI1.XI0.XI1<2>.XI7<1>.NET_003
+ XI1.XI0.XI1<2>.XI7<1>.NET_001 XI1.XI0.XI1<2>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_24 XI1.XI0.XI1<2>.XI7<1>.NET_004
+ XI1.XI0.XI1<2>.XI7<1>.NET_000 XI1.XI0.XI1<2>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<1>.NET_005
+ XI1.XI0.XI1<2>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<1>.NET_003
+ XI1.XI0.XI1<2>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_89_4 REG_DATA_2<1> XI1.XI0.XI1<2>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<1>.MM_i_55 XI1.XI0.XI1<2>.XI7<1>.NET_001
+ XI1.XI0.XI1<2>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_61 XI1.XI0.XI1<2>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_66 XI1.XI0.XI1<2>.XI7<1>.NET_003
+ XI1.XI0.XI1<2>.XI7<1>.NET_000 XI1.XI0.XI1<2>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_72 XI1.XI0.XI1<2>.XI7<1>.NET_007
+ XI1.XI0.XI1<2>.XI7<1>.NET_001 XI1.XI0.XI1<2>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<1>.NET_005
+ XI1.XI0.XI1<2>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<1>.NET_003
+ XI1.XI0.XI1<2>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_41_11 REG_DATA_2<0> XI1.XI0.XI1<2>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<0>.MM_i_7 XI1.XI0.XI1<2>.XI7<0>.NET_001
+ XI1.XI0.XI1<2>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_13 XI1.XI0.XI1<2>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_18 XI1.XI0.XI1<2>.XI7<0>.NET_003
+ XI1.XI0.XI1<2>.XI7<0>.NET_001 XI1.XI0.XI1<2>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_24 XI1.XI0.XI1<2>.XI7<0>.NET_004
+ XI1.XI0.XI1<2>.XI7<0>.NET_000 XI1.XI0.XI1<2>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<0>.NET_005
+ XI1.XI0.XI1<2>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<0>.NET_003
+ XI1.XI0.XI1<2>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_89_4 REG_DATA_2<0> XI1.XI0.XI1<2>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<0>.MM_i_55 XI1.XI0.XI1<2>.XI7<0>.NET_001
+ XI1.XI0.XI1<2>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_61 XI1.XI0.XI1<2>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_66 XI1.XI0.XI1<2>.XI7<0>.NET_003
+ XI1.XI0.XI1<2>.XI7<0>.NET_000 XI1.XI0.XI1<2>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_72 XI1.XI0.XI1<2>.XI7<0>.NET_007
+ XI1.XI0.XI1<2>.XI7<0>.NET_001 XI1.XI0.XI1<2>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<0>.NET_005
+ XI1.XI0.XI1<2>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<0>.NET_003
+ XI1.XI0.XI1<2>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_41_11 REG_DATA_2<7> XI1.XI0.XI1<2>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<7>.MM_i_7 XI1.XI0.XI1<2>.XI7<7>.NET_001
+ XI1.XI0.XI1<2>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_13 XI1.XI0.XI1<2>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_18 XI1.XI0.XI1<2>.XI7<7>.NET_003
+ XI1.XI0.XI1<2>.XI7<7>.NET_001 XI1.XI0.XI1<2>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_24 XI1.XI0.XI1<2>.XI7<7>.NET_004
+ XI1.XI0.XI1<2>.XI7<7>.NET_000 XI1.XI0.XI1<2>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<7>.NET_005
+ XI1.XI0.XI1<2>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<7>.NET_003
+ XI1.XI0.XI1<2>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_89_4 REG_DATA_2<7> XI1.XI0.XI1<2>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<7>.MM_i_55 XI1.XI0.XI1<2>.XI7<7>.NET_001
+ XI1.XI0.XI1<2>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_61 XI1.XI0.XI1<2>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_66 XI1.XI0.XI1<2>.XI7<7>.NET_003
+ XI1.XI0.XI1<2>.XI7<7>.NET_000 XI1.XI0.XI1<2>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_72 XI1.XI0.XI1<2>.XI7<7>.NET_007
+ XI1.XI0.XI1<2>.XI7<7>.NET_001 XI1.XI0.XI1<2>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<7>.NET_005
+ XI1.XI0.XI1<2>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<7>.NET_003
+ XI1.XI0.XI1<2>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_41_11 REG_DATA_2<6> XI1.XI0.XI1<2>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<6>.MM_i_7 XI1.XI0.XI1<2>.XI7<6>.NET_001
+ XI1.XI0.XI1<2>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_13 XI1.XI0.XI1<2>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_18 XI1.XI0.XI1<2>.XI7<6>.NET_003
+ XI1.XI0.XI1<2>.XI7<6>.NET_001 XI1.XI0.XI1<2>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_24 XI1.XI0.XI1<2>.XI7<6>.NET_004
+ XI1.XI0.XI1<2>.XI7<6>.NET_000 XI1.XI0.XI1<2>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<6>.NET_005
+ XI1.XI0.XI1<2>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<6>.NET_003
+ XI1.XI0.XI1<2>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_89_4 REG_DATA_2<6> XI1.XI0.XI1<2>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<6>.MM_i_55 XI1.XI0.XI1<2>.XI7<6>.NET_001
+ XI1.XI0.XI1<2>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_61 XI1.XI0.XI1<2>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_66 XI1.XI0.XI1<2>.XI7<6>.NET_003
+ XI1.XI0.XI1<2>.XI7<6>.NET_000 XI1.XI0.XI1<2>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_72 XI1.XI0.XI1<2>.XI7<6>.NET_007
+ XI1.XI0.XI1<2>.XI7<6>.NET_001 XI1.XI0.XI1<2>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<6>.NET_005
+ XI1.XI0.XI1<2>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<6>.NET_003
+ XI1.XI0.XI1<2>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_41_11 REG_DATA_2<5> XI1.XI0.XI1<2>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<5>.MM_i_7 XI1.XI0.XI1<2>.XI7<5>.NET_001
+ XI1.XI0.XI1<2>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_13 XI1.XI0.XI1<2>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_18 XI1.XI0.XI1<2>.XI7<5>.NET_003
+ XI1.XI0.XI1<2>.XI7<5>.NET_001 XI1.XI0.XI1<2>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_24 XI1.XI0.XI1<2>.XI7<5>.NET_004
+ XI1.XI0.XI1<2>.XI7<5>.NET_000 XI1.XI0.XI1<2>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<5>.NET_005
+ XI1.XI0.XI1<2>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<5>.NET_003
+ XI1.XI0.XI1<2>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_89_4 REG_DATA_2<5> XI1.XI0.XI1<2>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<5>.MM_i_55 XI1.XI0.XI1<2>.XI7<5>.NET_001
+ XI1.XI0.XI1<2>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_61 XI1.XI0.XI1<2>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_66 XI1.XI0.XI1<2>.XI7<5>.NET_003
+ XI1.XI0.XI1<2>.XI7<5>.NET_000 XI1.XI0.XI1<2>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_72 XI1.XI0.XI1<2>.XI7<5>.NET_007
+ XI1.XI0.XI1<2>.XI7<5>.NET_001 XI1.XI0.XI1<2>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<5>.NET_005
+ XI1.XI0.XI1<2>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<5>.NET_003
+ XI1.XI0.XI1<2>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_41_11 REG_DATA_2<4> XI1.XI0.XI1<2>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<4>.MM_i_7 XI1.XI0.XI1<2>.XI7<4>.NET_001
+ XI1.XI0.XI1<2>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_13 XI1.XI0.XI1<2>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_18 XI1.XI0.XI1<2>.XI7<4>.NET_003
+ XI1.XI0.XI1<2>.XI7<4>.NET_001 XI1.XI0.XI1<2>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_24 XI1.XI0.XI1<2>.XI7<4>.NET_004
+ XI1.XI0.XI1<2>.XI7<4>.NET_000 XI1.XI0.XI1<2>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<4>.NET_005
+ XI1.XI0.XI1<2>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<4>.NET_003
+ XI1.XI0.XI1<2>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_89_4 REG_DATA_2<4> XI1.XI0.XI1<2>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<4>.MM_i_55 XI1.XI0.XI1<2>.XI7<4>.NET_001
+ XI1.XI0.XI1<2>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_61 XI1.XI0.XI1<2>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_66 XI1.XI0.XI1<2>.XI7<4>.NET_003
+ XI1.XI0.XI1<2>.XI7<4>.NET_000 XI1.XI0.XI1<2>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_72 XI1.XI0.XI1<2>.XI7<4>.NET_007
+ XI1.XI0.XI1<2>.XI7<4>.NET_001 XI1.XI0.XI1<2>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<4>.NET_005
+ XI1.XI0.XI1<2>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<4>.NET_003
+ XI1.XI0.XI1<2>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_41_11 REG_DATA_2<11> XI1.XI0.XI1<2>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<11>.MM_i_7 XI1.XI0.XI1<2>.XI7<11>.NET_001
+ XI1.XI0.XI1<2>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_13 XI1.XI0.XI1<2>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_18 XI1.XI0.XI1<2>.XI7<11>.NET_003
+ XI1.XI0.XI1<2>.XI7<11>.NET_001 XI1.XI0.XI1<2>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_24 XI1.XI0.XI1<2>.XI7<11>.NET_004
+ XI1.XI0.XI1<2>.XI7<11>.NET_000 XI1.XI0.XI1<2>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<11>.NET_005
+ XI1.XI0.XI1<2>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<11>.NET_003
+ XI1.XI0.XI1<2>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_89_4 REG_DATA_2<11> XI1.XI0.XI1<2>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<11>.MM_i_55 XI1.XI0.XI1<2>.XI7<11>.NET_001
+ XI1.XI0.XI1<2>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_61 XI1.XI0.XI1<2>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_66 XI1.XI0.XI1<2>.XI7<11>.NET_003
+ XI1.XI0.XI1<2>.XI7<11>.NET_000 XI1.XI0.XI1<2>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_72 XI1.XI0.XI1<2>.XI7<11>.NET_007
+ XI1.XI0.XI1<2>.XI7<11>.NET_001 XI1.XI0.XI1<2>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<11>.NET_005
+ XI1.XI0.XI1<2>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<11>.NET_003
+ XI1.XI0.XI1<2>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_41_11 REG_DATA_2<10> XI1.XI0.XI1<2>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<10>.MM_i_7 XI1.XI0.XI1<2>.XI7<10>.NET_001
+ XI1.XI0.XI1<2>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_13 XI1.XI0.XI1<2>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_18 XI1.XI0.XI1<2>.XI7<10>.NET_003
+ XI1.XI0.XI1<2>.XI7<10>.NET_001 XI1.XI0.XI1<2>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_24 XI1.XI0.XI1<2>.XI7<10>.NET_004
+ XI1.XI0.XI1<2>.XI7<10>.NET_000 XI1.XI0.XI1<2>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<10>.NET_005
+ XI1.XI0.XI1<2>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<10>.NET_003
+ XI1.XI0.XI1<2>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_89_4 REG_DATA_2<10> XI1.XI0.XI1<2>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<10>.MM_i_55 XI1.XI0.XI1<2>.XI7<10>.NET_001
+ XI1.XI0.XI1<2>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_61 XI1.XI0.XI1<2>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_66 XI1.XI0.XI1<2>.XI7<10>.NET_003
+ XI1.XI0.XI1<2>.XI7<10>.NET_000 XI1.XI0.XI1<2>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_72 XI1.XI0.XI1<2>.XI7<10>.NET_007
+ XI1.XI0.XI1<2>.XI7<10>.NET_001 XI1.XI0.XI1<2>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<10>.NET_005
+ XI1.XI0.XI1<2>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<10>.NET_003
+ XI1.XI0.XI1<2>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_41_11 REG_DATA_2<9> XI1.XI0.XI1<2>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<9>.MM_i_7 XI1.XI0.XI1<2>.XI7<9>.NET_001
+ XI1.XI0.XI1<2>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_13 XI1.XI0.XI1<2>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_18 XI1.XI0.XI1<2>.XI7<9>.NET_003
+ XI1.XI0.XI1<2>.XI7<9>.NET_001 XI1.XI0.XI1<2>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_24 XI1.XI0.XI1<2>.XI7<9>.NET_004
+ XI1.XI0.XI1<2>.XI7<9>.NET_000 XI1.XI0.XI1<2>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<9>.NET_005
+ XI1.XI0.XI1<2>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<9>.NET_003
+ XI1.XI0.XI1<2>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_89_4 REG_DATA_2<9> XI1.XI0.XI1<2>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<9>.MM_i_55 XI1.XI0.XI1<2>.XI7<9>.NET_001
+ XI1.XI0.XI1<2>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_61 XI1.XI0.XI1<2>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_66 XI1.XI0.XI1<2>.XI7<9>.NET_003
+ XI1.XI0.XI1<2>.XI7<9>.NET_000 XI1.XI0.XI1<2>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_72 XI1.XI0.XI1<2>.XI7<9>.NET_007
+ XI1.XI0.XI1<2>.XI7<9>.NET_001 XI1.XI0.XI1<2>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<9>.NET_005
+ XI1.XI0.XI1<2>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<9>.NET_003
+ XI1.XI0.XI1<2>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_41_11 REG_DATA_2<8> XI1.XI0.XI1<2>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<8>.MM_i_7 XI1.XI0.XI1<2>.XI7<8>.NET_001
+ XI1.XI0.XI1<2>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_13 XI1.XI0.XI1<2>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_18 XI1.XI0.XI1<2>.XI7<8>.NET_003
+ XI1.XI0.XI1<2>.XI7<8>.NET_001 XI1.XI0.XI1<2>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_24 XI1.XI0.XI1<2>.XI7<8>.NET_004
+ XI1.XI0.XI1<2>.XI7<8>.NET_000 XI1.XI0.XI1<2>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<8>.NET_005
+ XI1.XI0.XI1<2>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<8>.NET_003
+ XI1.XI0.XI1<2>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_89_4 REG_DATA_2<8> XI1.XI0.XI1<2>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<8>.MM_i_55 XI1.XI0.XI1<2>.XI7<8>.NET_001
+ XI1.XI0.XI1<2>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_61 XI1.XI0.XI1<2>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_66 XI1.XI0.XI1<2>.XI7<8>.NET_003
+ XI1.XI0.XI1<2>.XI7<8>.NET_000 XI1.XI0.XI1<2>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_72 XI1.XI0.XI1<2>.XI7<8>.NET_007
+ XI1.XI0.XI1<2>.XI7<8>.NET_001 XI1.XI0.XI1<2>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<8>.NET_005
+ XI1.XI0.XI1<2>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<8>.NET_003
+ XI1.XI0.XI1<2>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_41_11 REG_DATA_2<15> XI1.XI0.XI1<2>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<15>.MM_i_7 XI1.XI0.XI1<2>.XI7<15>.NET_001
+ XI1.XI0.XI1<2>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_13 XI1.XI0.XI1<2>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_18 XI1.XI0.XI1<2>.XI7<15>.NET_003
+ XI1.XI0.XI1<2>.XI7<15>.NET_001 XI1.XI0.XI1<2>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_24 XI1.XI0.XI1<2>.XI7<15>.NET_004
+ XI1.XI0.XI1<2>.XI7<15>.NET_000 XI1.XI0.XI1<2>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<15>.NET_005
+ XI1.XI0.XI1<2>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<15>.NET_003
+ XI1.XI0.XI1<2>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_89_4 REG_DATA_2<15> XI1.XI0.XI1<2>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<15>.MM_i_55 XI1.XI0.XI1<2>.XI7<15>.NET_001
+ XI1.XI0.XI1<2>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_61 XI1.XI0.XI1<2>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_66 XI1.XI0.XI1<2>.XI7<15>.NET_003
+ XI1.XI0.XI1<2>.XI7<15>.NET_000 XI1.XI0.XI1<2>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_72 XI1.XI0.XI1<2>.XI7<15>.NET_007
+ XI1.XI0.XI1<2>.XI7<15>.NET_001 XI1.XI0.XI1<2>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<15>.NET_005
+ XI1.XI0.XI1<2>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<15>.NET_003
+ XI1.XI0.XI1<2>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_41_11 REG_DATA_2<14> XI1.XI0.XI1<2>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<14>.MM_i_7 XI1.XI0.XI1<2>.XI7<14>.NET_001
+ XI1.XI0.XI1<2>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_13 XI1.XI0.XI1<2>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_18 XI1.XI0.XI1<2>.XI7<14>.NET_003
+ XI1.XI0.XI1<2>.XI7<14>.NET_001 XI1.XI0.XI1<2>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_24 XI1.XI0.XI1<2>.XI7<14>.NET_004
+ XI1.XI0.XI1<2>.XI7<14>.NET_000 XI1.XI0.XI1<2>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<14>.NET_005
+ XI1.XI0.XI1<2>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<14>.NET_003
+ XI1.XI0.XI1<2>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_89_4 REG_DATA_2<14> XI1.XI0.XI1<2>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<14>.MM_i_55 XI1.XI0.XI1<2>.XI7<14>.NET_001
+ XI1.XI0.XI1<2>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_61 XI1.XI0.XI1<2>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_66 XI1.XI0.XI1<2>.XI7<14>.NET_003
+ XI1.XI0.XI1<2>.XI7<14>.NET_000 XI1.XI0.XI1<2>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_72 XI1.XI0.XI1<2>.XI7<14>.NET_007
+ XI1.XI0.XI1<2>.XI7<14>.NET_001 XI1.XI0.XI1<2>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<14>.NET_005
+ XI1.XI0.XI1<2>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<14>.NET_003
+ XI1.XI0.XI1<2>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_41_11 REG_DATA_2<13> XI1.XI0.XI1<2>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<13>.MM_i_7 XI1.XI0.XI1<2>.XI7<13>.NET_001
+ XI1.XI0.XI1<2>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_13 XI1.XI0.XI1<2>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_18 XI1.XI0.XI1<2>.XI7<13>.NET_003
+ XI1.XI0.XI1<2>.XI7<13>.NET_001 XI1.XI0.XI1<2>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_24 XI1.XI0.XI1<2>.XI7<13>.NET_004
+ XI1.XI0.XI1<2>.XI7<13>.NET_000 XI1.XI0.XI1<2>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<13>.NET_005
+ XI1.XI0.XI1<2>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<13>.NET_003
+ XI1.XI0.XI1<2>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_89_4 REG_DATA_2<13> XI1.XI0.XI1<2>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<13>.MM_i_55 XI1.XI0.XI1<2>.XI7<13>.NET_001
+ XI1.XI0.XI1<2>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_61 XI1.XI0.XI1<2>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_66 XI1.XI0.XI1<2>.XI7<13>.NET_003
+ XI1.XI0.XI1<2>.XI7<13>.NET_000 XI1.XI0.XI1<2>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_72 XI1.XI0.XI1<2>.XI7<13>.NET_007
+ XI1.XI0.XI1<2>.XI7<13>.NET_001 XI1.XI0.XI1<2>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<13>.NET_005
+ XI1.XI0.XI1<2>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<13>.NET_003
+ XI1.XI0.XI1<2>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_41_11 REG_DATA_2<12> XI1.XI0.XI1<2>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<2>.XI7<12>.MM_i_7 XI1.XI0.XI1<2>.XI7<12>.NET_001
+ XI1.XI0.XI1<2>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_13 XI1.XI0.XI1<2>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_18 XI1.XI0.XI1<2>.XI7<12>.NET_003
+ XI1.XI0.XI1<2>.XI7<12>.NET_001 XI1.XI0.XI1<2>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_24 XI1.XI0.XI1<2>.XI7<12>.NET_004
+ XI1.XI0.XI1<2>.XI7<12>.NET_000 XI1.XI0.XI1<2>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<2>.XI7<12>.NET_005
+ XI1.XI0.XI1<2>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<2>.XI7<12>.NET_003
+ XI1.XI0.XI1<2>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<2>
+ XI1.XI0.XI1<2>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_89_4 REG_DATA_2<12> XI1.XI0.XI1<2>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<2>.XI7<12>.MM_i_55 XI1.XI0.XI1<2>.XI7<12>.NET_001
+ XI1.XI0.XI1<2>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_61 XI1.XI0.XI1<2>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_66 XI1.XI0.XI1<2>.XI7<12>.NET_003
+ XI1.XI0.XI1<2>.XI7<12>.NET_000 XI1.XI0.XI1<2>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_72 XI1.XI0.XI1<2>.XI7<12>.NET_007
+ XI1.XI0.XI1<2>.XI7<12>.NET_001 XI1.XI0.XI1<2>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<2>.XI7<12>.NET_005
+ XI1.XI0.XI1<2>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<2>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<2>.XI7<12>.NET_003
+ XI1.XI0.XI1<2>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_41_11 REG_DATA_1<3> XI1.XI0.XI1<1>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<3>.MM_i_7 XI1.XI0.XI1<1>.XI7<3>.NET_001
+ XI1.XI0.XI1<1>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_13 XI1.XI0.XI1<1>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_18 XI1.XI0.XI1<1>.XI7<3>.NET_003
+ XI1.XI0.XI1<1>.XI7<3>.NET_001 XI1.XI0.XI1<1>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_24 XI1.XI0.XI1<1>.XI7<3>.NET_004
+ XI1.XI0.XI1<1>.XI7<3>.NET_000 XI1.XI0.XI1<1>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<3>.NET_005
+ XI1.XI0.XI1<1>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<3>.NET_003
+ XI1.XI0.XI1<1>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_89_4 REG_DATA_1<3> XI1.XI0.XI1<1>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<3>.MM_i_55 XI1.XI0.XI1<1>.XI7<3>.NET_001
+ XI1.XI0.XI1<1>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_61 XI1.XI0.XI1<1>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_66 XI1.XI0.XI1<1>.XI7<3>.NET_003
+ XI1.XI0.XI1<1>.XI7<3>.NET_000 XI1.XI0.XI1<1>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_72 XI1.XI0.XI1<1>.XI7<3>.NET_007
+ XI1.XI0.XI1<1>.XI7<3>.NET_001 XI1.XI0.XI1<1>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<3>.NET_005
+ XI1.XI0.XI1<1>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<3>.NET_003
+ XI1.XI0.XI1<1>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_41_11 REG_DATA_1<2> XI1.XI0.XI1<1>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<2>.MM_i_7 XI1.XI0.XI1<1>.XI7<2>.NET_001
+ XI1.XI0.XI1<1>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_13 XI1.XI0.XI1<1>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_18 XI1.XI0.XI1<1>.XI7<2>.NET_003
+ XI1.XI0.XI1<1>.XI7<2>.NET_001 XI1.XI0.XI1<1>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_24 XI1.XI0.XI1<1>.XI7<2>.NET_004
+ XI1.XI0.XI1<1>.XI7<2>.NET_000 XI1.XI0.XI1<1>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<2>.NET_005
+ XI1.XI0.XI1<1>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<2>.NET_003
+ XI1.XI0.XI1<1>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_89_4 REG_DATA_1<2> XI1.XI0.XI1<1>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<2>.MM_i_55 XI1.XI0.XI1<1>.XI7<2>.NET_001
+ XI1.XI0.XI1<1>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_61 XI1.XI0.XI1<1>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_66 XI1.XI0.XI1<1>.XI7<2>.NET_003
+ XI1.XI0.XI1<1>.XI7<2>.NET_000 XI1.XI0.XI1<1>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_72 XI1.XI0.XI1<1>.XI7<2>.NET_007
+ XI1.XI0.XI1<1>.XI7<2>.NET_001 XI1.XI0.XI1<1>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<2>.NET_005
+ XI1.XI0.XI1<1>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<2>.NET_003
+ XI1.XI0.XI1<1>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_41_11 REG_DATA_1<1> XI1.XI0.XI1<1>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<1>.MM_i_7 XI1.XI0.XI1<1>.XI7<1>.NET_001
+ XI1.XI0.XI1<1>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_13 XI1.XI0.XI1<1>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_18 XI1.XI0.XI1<1>.XI7<1>.NET_003
+ XI1.XI0.XI1<1>.XI7<1>.NET_001 XI1.XI0.XI1<1>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_24 XI1.XI0.XI1<1>.XI7<1>.NET_004
+ XI1.XI0.XI1<1>.XI7<1>.NET_000 XI1.XI0.XI1<1>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<1>.NET_005
+ XI1.XI0.XI1<1>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<1>.NET_003
+ XI1.XI0.XI1<1>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_89_4 REG_DATA_1<1> XI1.XI0.XI1<1>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<1>.MM_i_55 XI1.XI0.XI1<1>.XI7<1>.NET_001
+ XI1.XI0.XI1<1>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_61 XI1.XI0.XI1<1>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_66 XI1.XI0.XI1<1>.XI7<1>.NET_003
+ XI1.XI0.XI1<1>.XI7<1>.NET_000 XI1.XI0.XI1<1>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_72 XI1.XI0.XI1<1>.XI7<1>.NET_007
+ XI1.XI0.XI1<1>.XI7<1>.NET_001 XI1.XI0.XI1<1>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<1>.NET_005
+ XI1.XI0.XI1<1>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<1>.NET_003
+ XI1.XI0.XI1<1>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_41_11 REG_DATA_1<0> XI1.XI0.XI1<1>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<0>.MM_i_7 XI1.XI0.XI1<1>.XI7<0>.NET_001
+ XI1.XI0.XI1<1>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_13 XI1.XI0.XI1<1>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_18 XI1.XI0.XI1<1>.XI7<0>.NET_003
+ XI1.XI0.XI1<1>.XI7<0>.NET_001 XI1.XI0.XI1<1>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_24 XI1.XI0.XI1<1>.XI7<0>.NET_004
+ XI1.XI0.XI1<1>.XI7<0>.NET_000 XI1.XI0.XI1<1>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<0>.NET_005
+ XI1.XI0.XI1<1>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<0>.NET_003
+ XI1.XI0.XI1<1>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_89_4 REG_DATA_1<0> XI1.XI0.XI1<1>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<0>.MM_i_55 XI1.XI0.XI1<1>.XI7<0>.NET_001
+ XI1.XI0.XI1<1>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_61 XI1.XI0.XI1<1>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_66 XI1.XI0.XI1<1>.XI7<0>.NET_003
+ XI1.XI0.XI1<1>.XI7<0>.NET_000 XI1.XI0.XI1<1>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_72 XI1.XI0.XI1<1>.XI7<0>.NET_007
+ XI1.XI0.XI1<1>.XI7<0>.NET_001 XI1.XI0.XI1<1>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<0>.NET_005
+ XI1.XI0.XI1<1>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<0>.NET_003
+ XI1.XI0.XI1<1>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_41_11 REG_DATA_1<7> XI1.XI0.XI1<1>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<7>.MM_i_7 XI1.XI0.XI1<1>.XI7<7>.NET_001
+ XI1.XI0.XI1<1>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_13 XI1.XI0.XI1<1>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_18 XI1.XI0.XI1<1>.XI7<7>.NET_003
+ XI1.XI0.XI1<1>.XI7<7>.NET_001 XI1.XI0.XI1<1>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_24 XI1.XI0.XI1<1>.XI7<7>.NET_004
+ XI1.XI0.XI1<1>.XI7<7>.NET_000 XI1.XI0.XI1<1>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<7>.NET_005
+ XI1.XI0.XI1<1>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<7>.NET_003
+ XI1.XI0.XI1<1>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_89_4 REG_DATA_1<7> XI1.XI0.XI1<1>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<7>.MM_i_55 XI1.XI0.XI1<1>.XI7<7>.NET_001
+ XI1.XI0.XI1<1>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_61 XI1.XI0.XI1<1>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_66 XI1.XI0.XI1<1>.XI7<7>.NET_003
+ XI1.XI0.XI1<1>.XI7<7>.NET_000 XI1.XI0.XI1<1>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_72 XI1.XI0.XI1<1>.XI7<7>.NET_007
+ XI1.XI0.XI1<1>.XI7<7>.NET_001 XI1.XI0.XI1<1>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<7>.NET_005
+ XI1.XI0.XI1<1>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<7>.NET_003
+ XI1.XI0.XI1<1>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_41_11 REG_DATA_1<6> XI1.XI0.XI1<1>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<6>.MM_i_7 XI1.XI0.XI1<1>.XI7<6>.NET_001
+ XI1.XI0.XI1<1>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_13 XI1.XI0.XI1<1>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_18 XI1.XI0.XI1<1>.XI7<6>.NET_003
+ XI1.XI0.XI1<1>.XI7<6>.NET_001 XI1.XI0.XI1<1>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_24 XI1.XI0.XI1<1>.XI7<6>.NET_004
+ XI1.XI0.XI1<1>.XI7<6>.NET_000 XI1.XI0.XI1<1>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<6>.NET_005
+ XI1.XI0.XI1<1>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<6>.NET_003
+ XI1.XI0.XI1<1>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_89_4 REG_DATA_1<6> XI1.XI0.XI1<1>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<6>.MM_i_55 XI1.XI0.XI1<1>.XI7<6>.NET_001
+ XI1.XI0.XI1<1>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_61 XI1.XI0.XI1<1>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_66 XI1.XI0.XI1<1>.XI7<6>.NET_003
+ XI1.XI0.XI1<1>.XI7<6>.NET_000 XI1.XI0.XI1<1>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_72 XI1.XI0.XI1<1>.XI7<6>.NET_007
+ XI1.XI0.XI1<1>.XI7<6>.NET_001 XI1.XI0.XI1<1>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<6>.NET_005
+ XI1.XI0.XI1<1>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<6>.NET_003
+ XI1.XI0.XI1<1>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_41_11 REG_DATA_1<5> XI1.XI0.XI1<1>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<5>.MM_i_7 XI1.XI0.XI1<1>.XI7<5>.NET_001
+ XI1.XI0.XI1<1>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_13 XI1.XI0.XI1<1>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_18 XI1.XI0.XI1<1>.XI7<5>.NET_003
+ XI1.XI0.XI1<1>.XI7<5>.NET_001 XI1.XI0.XI1<1>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_24 XI1.XI0.XI1<1>.XI7<5>.NET_004
+ XI1.XI0.XI1<1>.XI7<5>.NET_000 XI1.XI0.XI1<1>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<5>.NET_005
+ XI1.XI0.XI1<1>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<5>.NET_003
+ XI1.XI0.XI1<1>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_89_4 REG_DATA_1<5> XI1.XI0.XI1<1>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<5>.MM_i_55 XI1.XI0.XI1<1>.XI7<5>.NET_001
+ XI1.XI0.XI1<1>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_61 XI1.XI0.XI1<1>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_66 XI1.XI0.XI1<1>.XI7<5>.NET_003
+ XI1.XI0.XI1<1>.XI7<5>.NET_000 XI1.XI0.XI1<1>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_72 XI1.XI0.XI1<1>.XI7<5>.NET_007
+ XI1.XI0.XI1<1>.XI7<5>.NET_001 XI1.XI0.XI1<1>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<5>.NET_005
+ XI1.XI0.XI1<1>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<5>.NET_003
+ XI1.XI0.XI1<1>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_41_11 REG_DATA_1<4> XI1.XI0.XI1<1>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<4>.MM_i_7 XI1.XI0.XI1<1>.XI7<4>.NET_001
+ XI1.XI0.XI1<1>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_13 XI1.XI0.XI1<1>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_18 XI1.XI0.XI1<1>.XI7<4>.NET_003
+ XI1.XI0.XI1<1>.XI7<4>.NET_001 XI1.XI0.XI1<1>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_24 XI1.XI0.XI1<1>.XI7<4>.NET_004
+ XI1.XI0.XI1<1>.XI7<4>.NET_000 XI1.XI0.XI1<1>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<4>.NET_005
+ XI1.XI0.XI1<1>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<4>.NET_003
+ XI1.XI0.XI1<1>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_89_4 REG_DATA_1<4> XI1.XI0.XI1<1>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<4>.MM_i_55 XI1.XI0.XI1<1>.XI7<4>.NET_001
+ XI1.XI0.XI1<1>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_61 XI1.XI0.XI1<1>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_66 XI1.XI0.XI1<1>.XI7<4>.NET_003
+ XI1.XI0.XI1<1>.XI7<4>.NET_000 XI1.XI0.XI1<1>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_72 XI1.XI0.XI1<1>.XI7<4>.NET_007
+ XI1.XI0.XI1<1>.XI7<4>.NET_001 XI1.XI0.XI1<1>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<4>.NET_005
+ XI1.XI0.XI1<1>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<4>.NET_003
+ XI1.XI0.XI1<1>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_41_11 REG_DATA_1<11> XI1.XI0.XI1<1>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<11>.MM_i_7 XI1.XI0.XI1<1>.XI7<11>.NET_001
+ XI1.XI0.XI1<1>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_13 XI1.XI0.XI1<1>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_18 XI1.XI0.XI1<1>.XI7<11>.NET_003
+ XI1.XI0.XI1<1>.XI7<11>.NET_001 XI1.XI0.XI1<1>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_24 XI1.XI0.XI1<1>.XI7<11>.NET_004
+ XI1.XI0.XI1<1>.XI7<11>.NET_000 XI1.XI0.XI1<1>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<11>.NET_005
+ XI1.XI0.XI1<1>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<11>.NET_003
+ XI1.XI0.XI1<1>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_89_4 REG_DATA_1<11> XI1.XI0.XI1<1>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<11>.MM_i_55 XI1.XI0.XI1<1>.XI7<11>.NET_001
+ XI1.XI0.XI1<1>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_61 XI1.XI0.XI1<1>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_66 XI1.XI0.XI1<1>.XI7<11>.NET_003
+ XI1.XI0.XI1<1>.XI7<11>.NET_000 XI1.XI0.XI1<1>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_72 XI1.XI0.XI1<1>.XI7<11>.NET_007
+ XI1.XI0.XI1<1>.XI7<11>.NET_001 XI1.XI0.XI1<1>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<11>.NET_005
+ XI1.XI0.XI1<1>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<11>.NET_003
+ XI1.XI0.XI1<1>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_41_11 REG_DATA_1<10> XI1.XI0.XI1<1>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<10>.MM_i_7 XI1.XI0.XI1<1>.XI7<10>.NET_001
+ XI1.XI0.XI1<1>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_13 XI1.XI0.XI1<1>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_18 XI1.XI0.XI1<1>.XI7<10>.NET_003
+ XI1.XI0.XI1<1>.XI7<10>.NET_001 XI1.XI0.XI1<1>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_24 XI1.XI0.XI1<1>.XI7<10>.NET_004
+ XI1.XI0.XI1<1>.XI7<10>.NET_000 XI1.XI0.XI1<1>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<10>.NET_005
+ XI1.XI0.XI1<1>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<10>.NET_003
+ XI1.XI0.XI1<1>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_89_4 REG_DATA_1<10> XI1.XI0.XI1<1>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<10>.MM_i_55 XI1.XI0.XI1<1>.XI7<10>.NET_001
+ XI1.XI0.XI1<1>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_61 XI1.XI0.XI1<1>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_66 XI1.XI0.XI1<1>.XI7<10>.NET_003
+ XI1.XI0.XI1<1>.XI7<10>.NET_000 XI1.XI0.XI1<1>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_72 XI1.XI0.XI1<1>.XI7<10>.NET_007
+ XI1.XI0.XI1<1>.XI7<10>.NET_001 XI1.XI0.XI1<1>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<10>.NET_005
+ XI1.XI0.XI1<1>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<10>.NET_003
+ XI1.XI0.XI1<1>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_41_11 REG_DATA_1<9> XI1.XI0.XI1<1>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<9>.MM_i_7 XI1.XI0.XI1<1>.XI7<9>.NET_001
+ XI1.XI0.XI1<1>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_13 XI1.XI0.XI1<1>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_18 XI1.XI0.XI1<1>.XI7<9>.NET_003
+ XI1.XI0.XI1<1>.XI7<9>.NET_001 XI1.XI0.XI1<1>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_24 XI1.XI0.XI1<1>.XI7<9>.NET_004
+ XI1.XI0.XI1<1>.XI7<9>.NET_000 XI1.XI0.XI1<1>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<9>.NET_005
+ XI1.XI0.XI1<1>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<9>.NET_003
+ XI1.XI0.XI1<1>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_89_4 REG_DATA_1<9> XI1.XI0.XI1<1>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<9>.MM_i_55 XI1.XI0.XI1<1>.XI7<9>.NET_001
+ XI1.XI0.XI1<1>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_61 XI1.XI0.XI1<1>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_66 XI1.XI0.XI1<1>.XI7<9>.NET_003
+ XI1.XI0.XI1<1>.XI7<9>.NET_000 XI1.XI0.XI1<1>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_72 XI1.XI0.XI1<1>.XI7<9>.NET_007
+ XI1.XI0.XI1<1>.XI7<9>.NET_001 XI1.XI0.XI1<1>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<9>.NET_005
+ XI1.XI0.XI1<1>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<9>.NET_003
+ XI1.XI0.XI1<1>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_41_11 REG_DATA_1<8> XI1.XI0.XI1<1>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<8>.MM_i_7 XI1.XI0.XI1<1>.XI7<8>.NET_001
+ XI1.XI0.XI1<1>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_13 XI1.XI0.XI1<1>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_18 XI1.XI0.XI1<1>.XI7<8>.NET_003
+ XI1.XI0.XI1<1>.XI7<8>.NET_001 XI1.XI0.XI1<1>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_24 XI1.XI0.XI1<1>.XI7<8>.NET_004
+ XI1.XI0.XI1<1>.XI7<8>.NET_000 XI1.XI0.XI1<1>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<8>.NET_005
+ XI1.XI0.XI1<1>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<8>.NET_003
+ XI1.XI0.XI1<1>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_89_4 REG_DATA_1<8> XI1.XI0.XI1<1>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<8>.MM_i_55 XI1.XI0.XI1<1>.XI7<8>.NET_001
+ XI1.XI0.XI1<1>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_61 XI1.XI0.XI1<1>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_66 XI1.XI0.XI1<1>.XI7<8>.NET_003
+ XI1.XI0.XI1<1>.XI7<8>.NET_000 XI1.XI0.XI1<1>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_72 XI1.XI0.XI1<1>.XI7<8>.NET_007
+ XI1.XI0.XI1<1>.XI7<8>.NET_001 XI1.XI0.XI1<1>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<8>.NET_005
+ XI1.XI0.XI1<1>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<8>.NET_003
+ XI1.XI0.XI1<1>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_41_11 REG_DATA_1<15> XI1.XI0.XI1<1>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<15>.MM_i_7 XI1.XI0.XI1<1>.XI7<15>.NET_001
+ XI1.XI0.XI1<1>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_13 XI1.XI0.XI1<1>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_18 XI1.XI0.XI1<1>.XI7<15>.NET_003
+ XI1.XI0.XI1<1>.XI7<15>.NET_001 XI1.XI0.XI1<1>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_24 XI1.XI0.XI1<1>.XI7<15>.NET_004
+ XI1.XI0.XI1<1>.XI7<15>.NET_000 XI1.XI0.XI1<1>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<15>.NET_005
+ XI1.XI0.XI1<1>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<15>.NET_003
+ XI1.XI0.XI1<1>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_89_4 REG_DATA_1<15> XI1.XI0.XI1<1>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<15>.MM_i_55 XI1.XI0.XI1<1>.XI7<15>.NET_001
+ XI1.XI0.XI1<1>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_61 XI1.XI0.XI1<1>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_66 XI1.XI0.XI1<1>.XI7<15>.NET_003
+ XI1.XI0.XI1<1>.XI7<15>.NET_000 XI1.XI0.XI1<1>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_72 XI1.XI0.XI1<1>.XI7<15>.NET_007
+ XI1.XI0.XI1<1>.XI7<15>.NET_001 XI1.XI0.XI1<1>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<15>.NET_005
+ XI1.XI0.XI1<1>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<15>.NET_003
+ XI1.XI0.XI1<1>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_41_11 REG_DATA_1<14> XI1.XI0.XI1<1>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<14>.MM_i_7 XI1.XI0.XI1<1>.XI7<14>.NET_001
+ XI1.XI0.XI1<1>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_13 XI1.XI0.XI1<1>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_18 XI1.XI0.XI1<1>.XI7<14>.NET_003
+ XI1.XI0.XI1<1>.XI7<14>.NET_001 XI1.XI0.XI1<1>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_24 XI1.XI0.XI1<1>.XI7<14>.NET_004
+ XI1.XI0.XI1<1>.XI7<14>.NET_000 XI1.XI0.XI1<1>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<14>.NET_005
+ XI1.XI0.XI1<1>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<14>.NET_003
+ XI1.XI0.XI1<1>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_89_4 REG_DATA_1<14> XI1.XI0.XI1<1>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<14>.MM_i_55 XI1.XI0.XI1<1>.XI7<14>.NET_001
+ XI1.XI0.XI1<1>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_61 XI1.XI0.XI1<1>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_66 XI1.XI0.XI1<1>.XI7<14>.NET_003
+ XI1.XI0.XI1<1>.XI7<14>.NET_000 XI1.XI0.XI1<1>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_72 XI1.XI0.XI1<1>.XI7<14>.NET_007
+ XI1.XI0.XI1<1>.XI7<14>.NET_001 XI1.XI0.XI1<1>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<14>.NET_005
+ XI1.XI0.XI1<1>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<14>.NET_003
+ XI1.XI0.XI1<1>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_41_11 REG_DATA_1<13> XI1.XI0.XI1<1>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<13>.MM_i_7 XI1.XI0.XI1<1>.XI7<13>.NET_001
+ XI1.XI0.XI1<1>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_13 XI1.XI0.XI1<1>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_18 XI1.XI0.XI1<1>.XI7<13>.NET_003
+ XI1.XI0.XI1<1>.XI7<13>.NET_001 XI1.XI0.XI1<1>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_24 XI1.XI0.XI1<1>.XI7<13>.NET_004
+ XI1.XI0.XI1<1>.XI7<13>.NET_000 XI1.XI0.XI1<1>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<13>.NET_005
+ XI1.XI0.XI1<1>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<13>.NET_003
+ XI1.XI0.XI1<1>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_89_4 REG_DATA_1<13> XI1.XI0.XI1<1>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<13>.MM_i_55 XI1.XI0.XI1<1>.XI7<13>.NET_001
+ XI1.XI0.XI1<1>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_61 XI1.XI0.XI1<1>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_66 XI1.XI0.XI1<1>.XI7<13>.NET_003
+ XI1.XI0.XI1<1>.XI7<13>.NET_000 XI1.XI0.XI1<1>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_72 XI1.XI0.XI1<1>.XI7<13>.NET_007
+ XI1.XI0.XI1<1>.XI7<13>.NET_001 XI1.XI0.XI1<1>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<13>.NET_005
+ XI1.XI0.XI1<1>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<13>.NET_003
+ XI1.XI0.XI1<1>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_41_11 REG_DATA_1<12> XI1.XI0.XI1<1>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<1>.XI7<12>.MM_i_7 XI1.XI0.XI1<1>.XI7<12>.NET_001
+ XI1.XI0.XI1<1>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_13 XI1.XI0.XI1<1>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_18 XI1.XI0.XI1<1>.XI7<12>.NET_003
+ XI1.XI0.XI1<1>.XI7<12>.NET_001 XI1.XI0.XI1<1>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_24 XI1.XI0.XI1<1>.XI7<12>.NET_004
+ XI1.XI0.XI1<1>.XI7<12>.NET_000 XI1.XI0.XI1<1>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<1>.XI7<12>.NET_005
+ XI1.XI0.XI1<1>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<1>.XI7<12>.NET_003
+ XI1.XI0.XI1<1>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<1>
+ XI1.XI0.XI1<1>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_89_4 REG_DATA_1<12> XI1.XI0.XI1<1>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<1>.XI7<12>.MM_i_55 XI1.XI0.XI1<1>.XI7<12>.NET_001
+ XI1.XI0.XI1<1>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_61 XI1.XI0.XI1<1>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_66 XI1.XI0.XI1<1>.XI7<12>.NET_003
+ XI1.XI0.XI1<1>.XI7<12>.NET_000 XI1.XI0.XI1<1>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_72 XI1.XI0.XI1<1>.XI7<12>.NET_007
+ XI1.XI0.XI1<1>.XI7<12>.NET_001 XI1.XI0.XI1<1>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<1>.XI7<12>.NET_005
+ XI1.XI0.XI1<1>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<1>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<1>.XI7<12>.NET_003
+ XI1.XI0.XI1<1>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<3>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_41_11 REG_DATA_0<3> XI1.XI0.XI1<0>.XI7<3>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<3>.MM_i_7 XI1.XI0.XI1<0>.XI7<3>.NET_001
+ XI1.XI0.XI1<0>.XI7<3>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_13 XI1.XI0.XI1<0>.XI7<3>.NET_002 XI1.XI0.M_DATA<3>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_18 XI1.XI0.XI1<0>.XI7<3>.NET_003
+ XI1.XI0.XI1<0>.XI7<3>.NET_001 XI1.XI0.XI1<0>.XI7<3>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_24 XI1.XI0.XI1<0>.XI7<3>.NET_004
+ XI1.XI0.XI1<0>.XI7<3>.NET_000 XI1.XI0.XI1<0>.XI7<3>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<3>.NET_005
+ XI1.XI0.XI1<0>.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<3>.NET_003
+ XI1.XI0.XI1<0>.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<3>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_89_4 REG_DATA_0<3> XI1.XI0.XI1<0>.XI7<3>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<3>.MM_i_55 XI1.XI0.XI1<0>.XI7<3>.NET_001
+ XI1.XI0.XI1<0>.XI7<3>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_61 XI1.XI0.XI1<0>.XI7<3>.NET_006 XI1.XI0.M_DATA<3>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_66 XI1.XI0.XI1<0>.XI7<3>.NET_003
+ XI1.XI0.XI1<0>.XI7<3>.NET_000 XI1.XI0.XI1<0>.XI7<3>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_72 XI1.XI0.XI1<0>.XI7<3>.NET_007
+ XI1.XI0.XI1<0>.XI7<3>.NET_001 XI1.XI0.XI1<0>.XI7<3>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<3>.NET_005
+ XI1.XI0.XI1<0>.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<3>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<3>.NET_003
+ XI1.XI0.XI1<0>.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<2>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_41_11 REG_DATA_0<2> XI1.XI0.XI1<0>.XI7<2>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<2>.MM_i_7 XI1.XI0.XI1<0>.XI7<2>.NET_001
+ XI1.XI0.XI1<0>.XI7<2>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_13 XI1.XI0.XI1<0>.XI7<2>.NET_002 XI1.XI0.M_DATA<2>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_18 XI1.XI0.XI1<0>.XI7<2>.NET_003
+ XI1.XI0.XI1<0>.XI7<2>.NET_001 XI1.XI0.XI1<0>.XI7<2>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_24 XI1.XI0.XI1<0>.XI7<2>.NET_004
+ XI1.XI0.XI1<0>.XI7<2>.NET_000 XI1.XI0.XI1<0>.XI7<2>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<2>.NET_005
+ XI1.XI0.XI1<0>.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<2>.NET_003
+ XI1.XI0.XI1<0>.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<2>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_89_4 REG_DATA_0<2> XI1.XI0.XI1<0>.XI7<2>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<2>.MM_i_55 XI1.XI0.XI1<0>.XI7<2>.NET_001
+ XI1.XI0.XI1<0>.XI7<2>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_61 XI1.XI0.XI1<0>.XI7<2>.NET_006 XI1.XI0.M_DATA<2>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_66 XI1.XI0.XI1<0>.XI7<2>.NET_003
+ XI1.XI0.XI1<0>.XI7<2>.NET_000 XI1.XI0.XI1<0>.XI7<2>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_72 XI1.XI0.XI1<0>.XI7<2>.NET_007
+ XI1.XI0.XI1<0>.XI7<2>.NET_001 XI1.XI0.XI1<0>.XI7<2>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<2>.NET_005
+ XI1.XI0.XI1<0>.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<2>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<2>.NET_003
+ XI1.XI0.XI1<0>.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<1>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_41_11 REG_DATA_0<1> XI1.XI0.XI1<0>.XI7<1>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<1>.MM_i_7 XI1.XI0.XI1<0>.XI7<1>.NET_001
+ XI1.XI0.XI1<0>.XI7<1>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_13 XI1.XI0.XI1<0>.XI7<1>.NET_002 XI1.XI0.M_DATA<1>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_18 XI1.XI0.XI1<0>.XI7<1>.NET_003
+ XI1.XI0.XI1<0>.XI7<1>.NET_001 XI1.XI0.XI1<0>.XI7<1>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_24 XI1.XI0.XI1<0>.XI7<1>.NET_004
+ XI1.XI0.XI1<0>.XI7<1>.NET_000 XI1.XI0.XI1<0>.XI7<1>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<1>.NET_005
+ XI1.XI0.XI1<0>.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<1>.NET_003
+ XI1.XI0.XI1<0>.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<1>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_89_4 REG_DATA_0<1> XI1.XI0.XI1<0>.XI7<1>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<1>.MM_i_55 XI1.XI0.XI1<0>.XI7<1>.NET_001
+ XI1.XI0.XI1<0>.XI7<1>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_61 XI1.XI0.XI1<0>.XI7<1>.NET_006 XI1.XI0.M_DATA<1>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_66 XI1.XI0.XI1<0>.XI7<1>.NET_003
+ XI1.XI0.XI1<0>.XI7<1>.NET_000 XI1.XI0.XI1<0>.XI7<1>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_72 XI1.XI0.XI1<0>.XI7<1>.NET_007
+ XI1.XI0.XI1<0>.XI7<1>.NET_001 XI1.XI0.XI1<0>.XI7<1>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<1>.NET_005
+ XI1.XI0.XI1<0>.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<1>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<1>.NET_003
+ XI1.XI0.XI1<0>.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<0>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_41_11 REG_DATA_0<0> XI1.XI0.XI1<0>.XI7<0>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<0>.MM_i_7 XI1.XI0.XI1<0>.XI7<0>.NET_001
+ XI1.XI0.XI1<0>.XI7<0>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_13 XI1.XI0.XI1<0>.XI7<0>.NET_002 XI1.XI0.M_DATA<0>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_18 XI1.XI0.XI1<0>.XI7<0>.NET_003
+ XI1.XI0.XI1<0>.XI7<0>.NET_001 XI1.XI0.XI1<0>.XI7<0>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_24 XI1.XI0.XI1<0>.XI7<0>.NET_004
+ XI1.XI0.XI1<0>.XI7<0>.NET_000 XI1.XI0.XI1<0>.XI7<0>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<0>.NET_005
+ XI1.XI0.XI1<0>.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<0>.NET_003
+ XI1.XI0.XI1<0>.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<0>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_89_4 REG_DATA_0<0> XI1.XI0.XI1<0>.XI7<0>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<0>.MM_i_55 XI1.XI0.XI1<0>.XI7<0>.NET_001
+ XI1.XI0.XI1<0>.XI7<0>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_61 XI1.XI0.XI1<0>.XI7<0>.NET_006 XI1.XI0.M_DATA<0>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_66 XI1.XI0.XI1<0>.XI7<0>.NET_003
+ XI1.XI0.XI1<0>.XI7<0>.NET_000 XI1.XI0.XI1<0>.XI7<0>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_72 XI1.XI0.XI1<0>.XI7<0>.NET_007
+ XI1.XI0.XI1<0>.XI7<0>.NET_001 XI1.XI0.XI1<0>.XI7<0>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<0>.NET_005
+ XI1.XI0.XI1<0>.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<0>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<0>.NET_003
+ XI1.XI0.XI1<0>.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<7>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_41_11 REG_DATA_0<7> XI1.XI0.XI1<0>.XI7<7>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<7>.MM_i_7 XI1.XI0.XI1<0>.XI7<7>.NET_001
+ XI1.XI0.XI1<0>.XI7<7>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_13 XI1.XI0.XI1<0>.XI7<7>.NET_002 XI1.XI0.M_DATA<7>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_18 XI1.XI0.XI1<0>.XI7<7>.NET_003
+ XI1.XI0.XI1<0>.XI7<7>.NET_001 XI1.XI0.XI1<0>.XI7<7>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_24 XI1.XI0.XI1<0>.XI7<7>.NET_004
+ XI1.XI0.XI1<0>.XI7<7>.NET_000 XI1.XI0.XI1<0>.XI7<7>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<7>.NET_005
+ XI1.XI0.XI1<0>.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<7>.NET_003
+ XI1.XI0.XI1<0>.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<7>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_89_4 REG_DATA_0<7> XI1.XI0.XI1<0>.XI7<7>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<7>.MM_i_55 XI1.XI0.XI1<0>.XI7<7>.NET_001
+ XI1.XI0.XI1<0>.XI7<7>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_61 XI1.XI0.XI1<0>.XI7<7>.NET_006 XI1.XI0.M_DATA<7>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_66 XI1.XI0.XI1<0>.XI7<7>.NET_003
+ XI1.XI0.XI1<0>.XI7<7>.NET_000 XI1.XI0.XI1<0>.XI7<7>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_72 XI1.XI0.XI1<0>.XI7<7>.NET_007
+ XI1.XI0.XI1<0>.XI7<7>.NET_001 XI1.XI0.XI1<0>.XI7<7>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<7>.NET_005
+ XI1.XI0.XI1<0>.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<7>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<7>.NET_003
+ XI1.XI0.XI1<0>.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<6>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_41_11 REG_DATA_0<6> XI1.XI0.XI1<0>.XI7<6>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<6>.MM_i_7 XI1.XI0.XI1<0>.XI7<6>.NET_001
+ XI1.XI0.XI1<0>.XI7<6>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_13 XI1.XI0.XI1<0>.XI7<6>.NET_002 XI1.XI0.M_DATA<6>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_18 XI1.XI0.XI1<0>.XI7<6>.NET_003
+ XI1.XI0.XI1<0>.XI7<6>.NET_001 XI1.XI0.XI1<0>.XI7<6>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_24 XI1.XI0.XI1<0>.XI7<6>.NET_004
+ XI1.XI0.XI1<0>.XI7<6>.NET_000 XI1.XI0.XI1<0>.XI7<6>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<6>.NET_005
+ XI1.XI0.XI1<0>.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<6>.NET_003
+ XI1.XI0.XI1<0>.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<6>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_89_4 REG_DATA_0<6> XI1.XI0.XI1<0>.XI7<6>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<6>.MM_i_55 XI1.XI0.XI1<0>.XI7<6>.NET_001
+ XI1.XI0.XI1<0>.XI7<6>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_61 XI1.XI0.XI1<0>.XI7<6>.NET_006 XI1.XI0.M_DATA<6>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_66 XI1.XI0.XI1<0>.XI7<6>.NET_003
+ XI1.XI0.XI1<0>.XI7<6>.NET_000 XI1.XI0.XI1<0>.XI7<6>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_72 XI1.XI0.XI1<0>.XI7<6>.NET_007
+ XI1.XI0.XI1<0>.XI7<6>.NET_001 XI1.XI0.XI1<0>.XI7<6>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<6>.NET_005
+ XI1.XI0.XI1<0>.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<6>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<6>.NET_003
+ XI1.XI0.XI1<0>.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<5>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_41_11 REG_DATA_0<5> XI1.XI0.XI1<0>.XI7<5>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<5>.MM_i_7 XI1.XI0.XI1<0>.XI7<5>.NET_001
+ XI1.XI0.XI1<0>.XI7<5>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_13 XI1.XI0.XI1<0>.XI7<5>.NET_002 XI1.XI0.M_DATA<5>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_18 XI1.XI0.XI1<0>.XI7<5>.NET_003
+ XI1.XI0.XI1<0>.XI7<5>.NET_001 XI1.XI0.XI1<0>.XI7<5>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_24 XI1.XI0.XI1<0>.XI7<5>.NET_004
+ XI1.XI0.XI1<0>.XI7<5>.NET_000 XI1.XI0.XI1<0>.XI7<5>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<5>.NET_005
+ XI1.XI0.XI1<0>.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<5>.NET_003
+ XI1.XI0.XI1<0>.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<5>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_89_4 REG_DATA_0<5> XI1.XI0.XI1<0>.XI7<5>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<5>.MM_i_55 XI1.XI0.XI1<0>.XI7<5>.NET_001
+ XI1.XI0.XI1<0>.XI7<5>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_61 XI1.XI0.XI1<0>.XI7<5>.NET_006 XI1.XI0.M_DATA<5>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_66 XI1.XI0.XI1<0>.XI7<5>.NET_003
+ XI1.XI0.XI1<0>.XI7<5>.NET_000 XI1.XI0.XI1<0>.XI7<5>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_72 XI1.XI0.XI1<0>.XI7<5>.NET_007
+ XI1.XI0.XI1<0>.XI7<5>.NET_001 XI1.XI0.XI1<0>.XI7<5>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<5>.NET_005
+ XI1.XI0.XI1<0>.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<5>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<5>.NET_003
+ XI1.XI0.XI1<0>.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<4>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_41_11 REG_DATA_0<4> XI1.XI0.XI1<0>.XI7<4>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<4>.MM_i_7 XI1.XI0.XI1<0>.XI7<4>.NET_001
+ XI1.XI0.XI1<0>.XI7<4>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_13 XI1.XI0.XI1<0>.XI7<4>.NET_002 XI1.XI0.M_DATA<4>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_18 XI1.XI0.XI1<0>.XI7<4>.NET_003
+ XI1.XI0.XI1<0>.XI7<4>.NET_001 XI1.XI0.XI1<0>.XI7<4>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_24 XI1.XI0.XI1<0>.XI7<4>.NET_004
+ XI1.XI0.XI1<0>.XI7<4>.NET_000 XI1.XI0.XI1<0>.XI7<4>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<4>.NET_005
+ XI1.XI0.XI1<0>.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<4>.NET_003
+ XI1.XI0.XI1<0>.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<4>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_89_4 REG_DATA_0<4> XI1.XI0.XI1<0>.XI7<4>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<4>.MM_i_55 XI1.XI0.XI1<0>.XI7<4>.NET_001
+ XI1.XI0.XI1<0>.XI7<4>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_61 XI1.XI0.XI1<0>.XI7<4>.NET_006 XI1.XI0.M_DATA<4>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_66 XI1.XI0.XI1<0>.XI7<4>.NET_003
+ XI1.XI0.XI1<0>.XI7<4>.NET_000 XI1.XI0.XI1<0>.XI7<4>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_72 XI1.XI0.XI1<0>.XI7<4>.NET_007
+ XI1.XI0.XI1<0>.XI7<4>.NET_001 XI1.XI0.XI1<0>.XI7<4>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<4>.NET_005
+ XI1.XI0.XI1<0>.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<4>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<4>.NET_003
+ XI1.XI0.XI1<0>.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<11>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_41_11 REG_DATA_0<11> XI1.XI0.XI1<0>.XI7<11>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<11>.MM_i_7 XI1.XI0.XI1<0>.XI7<11>.NET_001
+ XI1.XI0.XI1<0>.XI7<11>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_13 XI1.XI0.XI1<0>.XI7<11>.NET_002
+ XI1.XI0.M_DATA<11> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_18 XI1.XI0.XI1<0>.XI7<11>.NET_003
+ XI1.XI0.XI1<0>.XI7<11>.NET_001 XI1.XI0.XI1<0>.XI7<11>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_24 XI1.XI0.XI1<0>.XI7<11>.NET_004
+ XI1.XI0.XI1<0>.XI7<11>.NET_000 XI1.XI0.XI1<0>.XI7<11>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<11>.NET_005
+ XI1.XI0.XI1<0>.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<11>.NET_003
+ XI1.XI0.XI1<0>.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<11>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_89_4 REG_DATA_0<11> XI1.XI0.XI1<0>.XI7<11>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<11>.MM_i_55 XI1.XI0.XI1<0>.XI7<11>.NET_001
+ XI1.XI0.XI1<0>.XI7<11>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_61 XI1.XI0.XI1<0>.XI7<11>.NET_006
+ XI1.XI0.M_DATA<11> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_66 XI1.XI0.XI1<0>.XI7<11>.NET_003
+ XI1.XI0.XI1<0>.XI7<11>.NET_000 XI1.XI0.XI1<0>.XI7<11>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_72 XI1.XI0.XI1<0>.XI7<11>.NET_007
+ XI1.XI0.XI1<0>.XI7<11>.NET_001 XI1.XI0.XI1<0>.XI7<11>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<11>.NET_005
+ XI1.XI0.XI1<0>.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<11>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<11>.NET_003
+ XI1.XI0.XI1<0>.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<10>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_41_11 REG_DATA_0<10> XI1.XI0.XI1<0>.XI7<10>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<10>.MM_i_7 XI1.XI0.XI1<0>.XI7<10>.NET_001
+ XI1.XI0.XI1<0>.XI7<10>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_13 XI1.XI0.XI1<0>.XI7<10>.NET_002
+ XI1.XI0.M_DATA<10> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_18 XI1.XI0.XI1<0>.XI7<10>.NET_003
+ XI1.XI0.XI1<0>.XI7<10>.NET_001 XI1.XI0.XI1<0>.XI7<10>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_24 XI1.XI0.XI1<0>.XI7<10>.NET_004
+ XI1.XI0.XI1<0>.XI7<10>.NET_000 XI1.XI0.XI1<0>.XI7<10>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<10>.NET_005
+ XI1.XI0.XI1<0>.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<10>.NET_003
+ XI1.XI0.XI1<0>.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<10>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_89_4 REG_DATA_0<10> XI1.XI0.XI1<0>.XI7<10>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<10>.MM_i_55 XI1.XI0.XI1<0>.XI7<10>.NET_001
+ XI1.XI0.XI1<0>.XI7<10>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_61 XI1.XI0.XI1<0>.XI7<10>.NET_006
+ XI1.XI0.M_DATA<10> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_66 XI1.XI0.XI1<0>.XI7<10>.NET_003
+ XI1.XI0.XI1<0>.XI7<10>.NET_000 XI1.XI0.XI1<0>.XI7<10>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_72 XI1.XI0.XI1<0>.XI7<10>.NET_007
+ XI1.XI0.XI1<0>.XI7<10>.NET_001 XI1.XI0.XI1<0>.XI7<10>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<10>.NET_005
+ XI1.XI0.XI1<0>.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<10>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<10>.NET_003
+ XI1.XI0.XI1<0>.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<9>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_41_11 REG_DATA_0<9> XI1.XI0.XI1<0>.XI7<9>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<9>.MM_i_7 XI1.XI0.XI1<0>.XI7<9>.NET_001
+ XI1.XI0.XI1<0>.XI7<9>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_13 XI1.XI0.XI1<0>.XI7<9>.NET_002 XI1.XI0.M_DATA<9>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_18 XI1.XI0.XI1<0>.XI7<9>.NET_003
+ XI1.XI0.XI1<0>.XI7<9>.NET_001 XI1.XI0.XI1<0>.XI7<9>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_24 XI1.XI0.XI1<0>.XI7<9>.NET_004
+ XI1.XI0.XI1<0>.XI7<9>.NET_000 XI1.XI0.XI1<0>.XI7<9>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<9>.NET_005
+ XI1.XI0.XI1<0>.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<9>.NET_003
+ XI1.XI0.XI1<0>.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<9>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_89_4 REG_DATA_0<9> XI1.XI0.XI1<0>.XI7<9>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<9>.MM_i_55 XI1.XI0.XI1<0>.XI7<9>.NET_001
+ XI1.XI0.XI1<0>.XI7<9>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_61 XI1.XI0.XI1<0>.XI7<9>.NET_006 XI1.XI0.M_DATA<9>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_66 XI1.XI0.XI1<0>.XI7<9>.NET_003
+ XI1.XI0.XI1<0>.XI7<9>.NET_000 XI1.XI0.XI1<0>.XI7<9>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_72 XI1.XI0.XI1<0>.XI7<9>.NET_007
+ XI1.XI0.XI1<0>.XI7<9>.NET_001 XI1.XI0.XI1<0>.XI7<9>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<9>.NET_005
+ XI1.XI0.XI1<0>.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<9>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<9>.NET_003
+ XI1.XI0.XI1<0>.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<8>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_41_11 REG_DATA_0<8> XI1.XI0.XI1<0>.XI7<8>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<8>.MM_i_7 XI1.XI0.XI1<0>.XI7<8>.NET_001
+ XI1.XI0.XI1<0>.XI7<8>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_13 XI1.XI0.XI1<0>.XI7<8>.NET_002 XI1.XI0.M_DATA<8>
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_18 XI1.XI0.XI1<0>.XI7<8>.NET_003
+ XI1.XI0.XI1<0>.XI7<8>.NET_001 XI1.XI0.XI1<0>.XI7<8>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_24 XI1.XI0.XI1<0>.XI7<8>.NET_004
+ XI1.XI0.XI1<0>.XI7<8>.NET_000 XI1.XI0.XI1<0>.XI7<8>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<8>.NET_005
+ XI1.XI0.XI1<0>.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<8>.NET_003
+ XI1.XI0.XI1<0>.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<8>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_89_4 REG_DATA_0<8> XI1.XI0.XI1<0>.XI7<8>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<8>.MM_i_55 XI1.XI0.XI1<0>.XI7<8>.NET_001
+ XI1.XI0.XI1<0>.XI7<8>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_61 XI1.XI0.XI1<0>.XI7<8>.NET_006 XI1.XI0.M_DATA<8>
+ VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07
+ PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_66 XI1.XI0.XI1<0>.XI7<8>.NET_003
+ XI1.XI0.XI1<0>.XI7<8>.NET_000 XI1.XI0.XI1<0>.XI7<8>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_72 XI1.XI0.XI1<0>.XI7<8>.NET_007
+ XI1.XI0.XI1<0>.XI7<8>.NET_001 XI1.XI0.XI1<0>.XI7<8>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<8>.NET_005
+ XI1.XI0.XI1<0>.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<8>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<8>.NET_003
+ XI1.XI0.XI1<0>.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<15>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_41_11 REG_DATA_0<15> XI1.XI0.XI1<0>.XI7<15>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<15>.MM_i_7 XI1.XI0.XI1<0>.XI7<15>.NET_001
+ XI1.XI0.XI1<0>.XI7<15>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_13 XI1.XI0.XI1<0>.XI7<15>.NET_002
+ XI1.XI0.M_DATA<15> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_18 XI1.XI0.XI1<0>.XI7<15>.NET_003
+ XI1.XI0.XI1<0>.XI7<15>.NET_001 XI1.XI0.XI1<0>.XI7<15>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_24 XI1.XI0.XI1<0>.XI7<15>.NET_004
+ XI1.XI0.XI1<0>.XI7<15>.NET_000 XI1.XI0.XI1<0>.XI7<15>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<15>.NET_005
+ XI1.XI0.XI1<0>.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<15>.NET_003
+ XI1.XI0.XI1<0>.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<15>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_89_4 REG_DATA_0<15> XI1.XI0.XI1<0>.XI7<15>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<15>.MM_i_55 XI1.XI0.XI1<0>.XI7<15>.NET_001
+ XI1.XI0.XI1<0>.XI7<15>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_61 XI1.XI0.XI1<0>.XI7<15>.NET_006
+ XI1.XI0.M_DATA<15> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_66 XI1.XI0.XI1<0>.XI7<15>.NET_003
+ XI1.XI0.XI1<0>.XI7<15>.NET_000 XI1.XI0.XI1<0>.XI7<15>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_72 XI1.XI0.XI1<0>.XI7<15>.NET_007
+ XI1.XI0.XI1<0>.XI7<15>.NET_001 XI1.XI0.XI1<0>.XI7<15>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<15>.NET_005
+ XI1.XI0.XI1<0>.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<15>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<15>.NET_003
+ XI1.XI0.XI1<0>.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<14>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_41_11 REG_DATA_0<14> XI1.XI0.XI1<0>.XI7<14>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<14>.MM_i_7 XI1.XI0.XI1<0>.XI7<14>.NET_001
+ XI1.XI0.XI1<0>.XI7<14>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_13 XI1.XI0.XI1<0>.XI7<14>.NET_002
+ XI1.XI0.M_DATA<14> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_18 XI1.XI0.XI1<0>.XI7<14>.NET_003
+ XI1.XI0.XI1<0>.XI7<14>.NET_001 XI1.XI0.XI1<0>.XI7<14>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_24 XI1.XI0.XI1<0>.XI7<14>.NET_004
+ XI1.XI0.XI1<0>.XI7<14>.NET_000 XI1.XI0.XI1<0>.XI7<14>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<14>.NET_005
+ XI1.XI0.XI1<0>.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<14>.NET_003
+ XI1.XI0.XI1<0>.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<14>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_89_4 REG_DATA_0<14> XI1.XI0.XI1<0>.XI7<14>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<14>.MM_i_55 XI1.XI0.XI1<0>.XI7<14>.NET_001
+ XI1.XI0.XI1<0>.XI7<14>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_61 XI1.XI0.XI1<0>.XI7<14>.NET_006
+ XI1.XI0.M_DATA<14> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_66 XI1.XI0.XI1<0>.XI7<14>.NET_003
+ XI1.XI0.XI1<0>.XI7<14>.NET_000 XI1.XI0.XI1<0>.XI7<14>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_72 XI1.XI0.XI1<0>.XI7<14>.NET_007
+ XI1.XI0.XI1<0>.XI7<14>.NET_001 XI1.XI0.XI1<0>.XI7<14>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<14>.NET_005
+ XI1.XI0.XI1<0>.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<14>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<14>.NET_003
+ XI1.XI0.XI1<0>.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<13>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_41_11 REG_DATA_0<13> XI1.XI0.XI1<0>.XI7<13>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<13>.MM_i_7 XI1.XI0.XI1<0>.XI7<13>.NET_001
+ XI1.XI0.XI1<0>.XI7<13>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_13 XI1.XI0.XI1<0>.XI7<13>.NET_002
+ XI1.XI0.M_DATA<13> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_18 XI1.XI0.XI1<0>.XI7<13>.NET_003
+ XI1.XI0.XI1<0>.XI7<13>.NET_001 XI1.XI0.XI1<0>.XI7<13>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_24 XI1.XI0.XI1<0>.XI7<13>.NET_004
+ XI1.XI0.XI1<0>.XI7<13>.NET_000 XI1.XI0.XI1<0>.XI7<13>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<13>.NET_005
+ XI1.XI0.XI1<0>.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<13>.NET_003
+ XI1.XI0.XI1<0>.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<13>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_89_4 REG_DATA_0<13> XI1.XI0.XI1<0>.XI7<13>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<13>.MM_i_55 XI1.XI0.XI1<0>.XI7<13>.NET_001
+ XI1.XI0.XI1<0>.XI7<13>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_61 XI1.XI0.XI1<0>.XI7<13>.NET_006
+ XI1.XI0.M_DATA<13> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_66 XI1.XI0.XI1<0>.XI7<13>.NET_003
+ XI1.XI0.XI1<0>.XI7<13>.NET_000 XI1.XI0.XI1<0>.XI7<13>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_72 XI1.XI0.XI1<0>.XI7<13>.NET_007
+ XI1.XI0.XI1<0>.XI7<13>.NET_001 XI1.XI0.XI1<0>.XI7<13>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<13>.NET_005
+ XI1.XI0.XI1<0>.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<13>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<13>.NET_003
+ XI1.XI0.XI1<0>.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_0 VSS! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<12>.NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.205e-14 PD=1.11e-06 PS=6.3e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_41_11 REG_DATA_0<12> XI1.XI0.XI1<0>.XI7<12>.NET_003
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI1<0>.XI7<12>.MM_i_7 XI1.XI0.XI1<0>.XI7<12>.NET_001
+ XI1.XI0.XI1<0>.XI7<12>.NET_000 VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_13 XI1.XI0.XI1<0>.XI7<12>.NET_002
+ XI1.XI0.M_DATA<12> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_18 XI1.XI0.XI1<0>.XI7<12>.NET_003
+ XI1.XI0.XI1<0>.XI7<12>.NET_001 XI1.XI0.XI1<0>.XI7<12>.NET_002 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_24 XI1.XI0.XI1<0>.XI7<12>.NET_004
+ XI1.XI0.XI1<0>.XI7<12>.NET_000 XI1.XI0.XI1<0>.XI7<12>.NET_003 VSS! NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_28 VSS! XI1.XI0.XI1<0>.XI7<12>.NET_005
+ XI1.XI0.XI1<0>.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_34 VSS! XI1.XI0.XI1<0>.XI7<12>.NET_003
+ XI1.XI0.XI1<0>.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_48 VDD! XI1.XI0.CK_EN<0>
+ XI1.XI0.XI1<0>.XI7<12>.NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_89_4 REG_DATA_0<12> XI1.XI0.XI1<0>.XI7<12>.NET_003
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI1<0>.XI7<12>.MM_i_55 XI1.XI0.XI1<0>.XI7<12>.NET_001
+ XI1.XI0.XI1<0>.XI7<12>.NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_61 XI1.XI0.XI1<0>.XI7<12>.NET_006
+ XI1.XI0.M_DATA<12> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_66 XI1.XI0.XI1<0>.XI7<12>.NET_003
+ XI1.XI0.XI1<0>.XI7<12>.NET_000 XI1.XI0.XI1<0>.XI7<12>.NET_006 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_72 XI1.XI0.XI1<0>.XI7<12>.NET_007
+ XI1.XI0.XI1<0>.XI7<12>.NET_001 XI1.XI0.XI1<0>.XI7<12>.NET_003 VDD! PMOS_VTL
+ L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_76 VDD! XI1.XI0.XI1<0>.XI7<12>.NET_005
+ XI1.XI0.XI1<0>.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI1<0>.XI7<12>.MM_i_82 VDD! XI1.XI0.XI1<0>.XI7<12>.NET_003
+ XI1.XI0.XI1<0>.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI16.MM_i_2 XI1.XI0.NET5 XI1.XI0.CK_EN<12> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI16.MM_i_1 VSS! XI1.XI0.CK_EN<11> XI1.XI0.NET5 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI16.MM_i_0 XI1.XI0.NET5 XI1.XI0.CK_EN<10> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI16.MM_i_5 XI1.XI0.XI16.NET_1 XI1.XI0.CK_EN<12> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI16.MM_i_4 XI1.XI0.XI16.NET_0 XI1.XI0.CK_EN<11> XI1.XI0.XI16.NET_1
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI1.XI0.XI16.MM_i_3 XI1.XI0.NET5 XI1.XI0.CK_EN<10> XI1.XI0.XI16.NET_0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI17.MM_i_2 XI1.XI0.NET13 XI1.XI0.CK_EN<7> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI17.MM_i_1 VSS! XI1.XI0.CK_EN<9> XI1.XI0.NET13 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI17.MM_i_0 XI1.XI0.NET13 XI1.XI0.CK_EN<8> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI17.MM_i_5 XI1.XI0.XI17.NET_1 XI1.XI0.CK_EN<7> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI17.MM_i_4 XI1.XI0.XI17.NET_0 XI1.XI0.CK_EN<9> XI1.XI0.XI17.NET_1 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI17.MM_i_3 XI1.XI0.NET13 XI1.XI0.CK_EN<8> XI1.XI0.XI17.NET_0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI15.MM_i_2 XI1.XI0.NET9 XI1.XI0.CK_EN<6> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI1.XI0.XI15.MM_i_1 VSS! XI1.XI0.CK_EN<5> XI1.XI0.NET9 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI1.XI0.XI15.MM_i_0 XI1.XI0.NET9 XI1.XI0.CK_EN<4> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI1.XI0.XI15.MM_i_5 XI1.XI0.XI15.NET_1 XI1.XI0.CK_EN<6> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI15.MM_i_4 XI1.XI0.XI15.NET_0 XI1.XI0.CK_EN<5> XI1.XI0.XI15.NET_1 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI15.MM_i_3 XI1.XI0.NET9 XI1.XI0.CK_EN<4> XI1.XI0.XI15.NET_0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI0.XI7<3>.MM_i_7 VSS! XI1.XI0.XI0.XI7<3>.NET_000
+ XI1.XI0.XI0.XI7<3>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<3>.MM_i_13 XI1.XI0.XI0.XI7<3>.NET_002 WR_DATA<3> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<3>.MM_i_18 XI1.XI0.XI0.XI7<3>.NET_003
+ XI1.XI0.XI0.XI7<3>.NET_000 XI1.XI0.XI0.XI7<3>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<3>.MM_i_24 XI1.XI0.XI0.XI7<3>.NET_004
+ XI1.XI0.XI0.XI7<3>.NET_001 XI1.XI0.XI0.XI7<3>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<3>.MM_i_29 VSS! XI1.XI0.XI0.XI7<3>.NET_005
+ XI1.XI0.XI0.XI7<3>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<3>.MM_i_35 VSS! XI1.XI0.XI0.XI7<3>.NET_003
+ XI1.XI0.XI0.XI7<3>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<3>.MM_i_42 XI1.XI0.M_DATA<3> XI1.XI0.XI0.XI7<3>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<3>.MM_i_0 XI1.XI0.XI0.XI7<3>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<3>.MM_i_55 VDD! XI1.XI0.XI0.XI7<3>.NET_000
+ XI1.XI0.XI0.XI7<3>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<3>.MM_i_62 XI1.XI0.XI0.XI7<3>.NET_006 WR_DATA<3> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<3>.MM_i_67 XI1.XI0.XI0.XI7<3>.NET_003
+ XI1.XI0.XI0.XI7<3>.NET_001 XI1.XI0.XI0.XI7<3>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<3>.MM_i_73 XI1.XI0.XI0.XI7<3>.NET_007
+ XI1.XI0.XI0.XI7<3>.NET_000 XI1.XI0.XI0.XI7<3>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<3>.MM_i_79 VDD! XI1.XI0.XI0.XI7<3>.NET_005
+ XI1.XI0.XI0.XI7<3>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<3>.MM_i_85 VDD! XI1.XI0.XI0.XI7<3>.NET_003
+ XI1.XI0.XI0.XI7<3>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<3>.MM_i_92 XI1.XI0.M_DATA<3> XI1.XI0.XI0.XI7<3>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<3>.MM_i_48 XI1.XI0.XI0.XI7<3>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<2>.MM_i_7 VSS! XI1.XI0.XI0.XI7<2>.NET_000
+ XI1.XI0.XI0.XI7<2>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<2>.MM_i_13 XI1.XI0.XI0.XI7<2>.NET_002 WR_DATA<2> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<2>.MM_i_18 XI1.XI0.XI0.XI7<2>.NET_003
+ XI1.XI0.XI0.XI7<2>.NET_000 XI1.XI0.XI0.XI7<2>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<2>.MM_i_24 XI1.XI0.XI0.XI7<2>.NET_004
+ XI1.XI0.XI0.XI7<2>.NET_001 XI1.XI0.XI0.XI7<2>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<2>.MM_i_29 VSS! XI1.XI0.XI0.XI7<2>.NET_005
+ XI1.XI0.XI0.XI7<2>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<2>.MM_i_35 VSS! XI1.XI0.XI0.XI7<2>.NET_003
+ XI1.XI0.XI0.XI7<2>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<2>.MM_i_42 XI1.XI0.M_DATA<2> XI1.XI0.XI0.XI7<2>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<2>.MM_i_0 XI1.XI0.XI0.XI7<2>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<2>.MM_i_55 VDD! XI1.XI0.XI0.XI7<2>.NET_000
+ XI1.XI0.XI0.XI7<2>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<2>.MM_i_62 XI1.XI0.XI0.XI7<2>.NET_006 WR_DATA<2> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<2>.MM_i_67 XI1.XI0.XI0.XI7<2>.NET_003
+ XI1.XI0.XI0.XI7<2>.NET_001 XI1.XI0.XI0.XI7<2>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<2>.MM_i_73 XI1.XI0.XI0.XI7<2>.NET_007
+ XI1.XI0.XI0.XI7<2>.NET_000 XI1.XI0.XI0.XI7<2>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<2>.MM_i_79 VDD! XI1.XI0.XI0.XI7<2>.NET_005
+ XI1.XI0.XI0.XI7<2>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<2>.MM_i_85 VDD! XI1.XI0.XI0.XI7<2>.NET_003
+ XI1.XI0.XI0.XI7<2>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<2>.MM_i_92 XI1.XI0.M_DATA<2> XI1.XI0.XI0.XI7<2>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<2>.MM_i_48 XI1.XI0.XI0.XI7<2>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<1>.MM_i_7 VSS! XI1.XI0.XI0.XI7<1>.NET_000
+ XI1.XI0.XI0.XI7<1>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<1>.MM_i_13 XI1.XI0.XI0.XI7<1>.NET_002 WR_DATA<1> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<1>.MM_i_18 XI1.XI0.XI0.XI7<1>.NET_003
+ XI1.XI0.XI0.XI7<1>.NET_000 XI1.XI0.XI0.XI7<1>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<1>.MM_i_24 XI1.XI0.XI0.XI7<1>.NET_004
+ XI1.XI0.XI0.XI7<1>.NET_001 XI1.XI0.XI0.XI7<1>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<1>.MM_i_29 VSS! XI1.XI0.XI0.XI7<1>.NET_005
+ XI1.XI0.XI0.XI7<1>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<1>.MM_i_35 VSS! XI1.XI0.XI0.XI7<1>.NET_003
+ XI1.XI0.XI0.XI7<1>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<1>.MM_i_42 XI1.XI0.M_DATA<1> XI1.XI0.XI0.XI7<1>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<1>.MM_i_0 XI1.XI0.XI0.XI7<1>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<1>.MM_i_55 VDD! XI1.XI0.XI0.XI7<1>.NET_000
+ XI1.XI0.XI0.XI7<1>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<1>.MM_i_62 XI1.XI0.XI0.XI7<1>.NET_006 WR_DATA<1> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<1>.MM_i_67 XI1.XI0.XI0.XI7<1>.NET_003
+ XI1.XI0.XI0.XI7<1>.NET_001 XI1.XI0.XI0.XI7<1>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<1>.MM_i_73 XI1.XI0.XI0.XI7<1>.NET_007
+ XI1.XI0.XI0.XI7<1>.NET_000 XI1.XI0.XI0.XI7<1>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<1>.MM_i_79 VDD! XI1.XI0.XI0.XI7<1>.NET_005
+ XI1.XI0.XI0.XI7<1>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<1>.MM_i_85 VDD! XI1.XI0.XI0.XI7<1>.NET_003
+ XI1.XI0.XI0.XI7<1>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<1>.MM_i_92 XI1.XI0.M_DATA<1> XI1.XI0.XI0.XI7<1>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<1>.MM_i_48 XI1.XI0.XI0.XI7<1>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<0>.MM_i_7 VSS! XI1.XI0.XI0.XI7<0>.NET_000
+ XI1.XI0.XI0.XI7<0>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<0>.MM_i_13 XI1.XI0.XI0.XI7<0>.NET_002 WR_DATA<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<0>.MM_i_18 XI1.XI0.XI0.XI7<0>.NET_003
+ XI1.XI0.XI0.XI7<0>.NET_000 XI1.XI0.XI0.XI7<0>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<0>.MM_i_24 XI1.XI0.XI0.XI7<0>.NET_004
+ XI1.XI0.XI0.XI7<0>.NET_001 XI1.XI0.XI0.XI7<0>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<0>.MM_i_29 VSS! XI1.XI0.XI0.XI7<0>.NET_005
+ XI1.XI0.XI0.XI7<0>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<0>.MM_i_35 VSS! XI1.XI0.XI0.XI7<0>.NET_003
+ XI1.XI0.XI0.XI7<0>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<0>.MM_i_42 XI1.XI0.M_DATA<0> XI1.XI0.XI0.XI7<0>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<0>.MM_i_0 XI1.XI0.XI0.XI7<0>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<0>.MM_i_55 VDD! XI1.XI0.XI0.XI7<0>.NET_000
+ XI1.XI0.XI0.XI7<0>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<0>.MM_i_62 XI1.XI0.XI0.XI7<0>.NET_006 WR_DATA<0> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<0>.MM_i_67 XI1.XI0.XI0.XI7<0>.NET_003
+ XI1.XI0.XI0.XI7<0>.NET_001 XI1.XI0.XI0.XI7<0>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<0>.MM_i_73 XI1.XI0.XI0.XI7<0>.NET_007
+ XI1.XI0.XI0.XI7<0>.NET_000 XI1.XI0.XI0.XI7<0>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<0>.MM_i_79 VDD! XI1.XI0.XI0.XI7<0>.NET_005
+ XI1.XI0.XI0.XI7<0>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<0>.MM_i_85 VDD! XI1.XI0.XI0.XI7<0>.NET_003
+ XI1.XI0.XI0.XI7<0>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<0>.MM_i_92 XI1.XI0.M_DATA<0> XI1.XI0.XI0.XI7<0>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<0>.MM_i_48 XI1.XI0.XI0.XI7<0>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<7>.MM_i_7 VSS! XI1.XI0.XI0.XI7<7>.NET_000
+ XI1.XI0.XI0.XI7<7>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<7>.MM_i_13 XI1.XI0.XI0.XI7<7>.NET_002 WR_DATA<7> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<7>.MM_i_18 XI1.XI0.XI0.XI7<7>.NET_003
+ XI1.XI0.XI0.XI7<7>.NET_000 XI1.XI0.XI0.XI7<7>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<7>.MM_i_24 XI1.XI0.XI0.XI7<7>.NET_004
+ XI1.XI0.XI0.XI7<7>.NET_001 XI1.XI0.XI0.XI7<7>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<7>.MM_i_29 VSS! XI1.XI0.XI0.XI7<7>.NET_005
+ XI1.XI0.XI0.XI7<7>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<7>.MM_i_35 VSS! XI1.XI0.XI0.XI7<7>.NET_003
+ XI1.XI0.XI0.XI7<7>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<7>.MM_i_42 XI1.XI0.M_DATA<7> XI1.XI0.XI0.XI7<7>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<7>.MM_i_0 XI1.XI0.XI0.XI7<7>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<7>.MM_i_55 VDD! XI1.XI0.XI0.XI7<7>.NET_000
+ XI1.XI0.XI0.XI7<7>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<7>.MM_i_62 XI1.XI0.XI0.XI7<7>.NET_006 WR_DATA<7> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<7>.MM_i_67 XI1.XI0.XI0.XI7<7>.NET_003
+ XI1.XI0.XI0.XI7<7>.NET_001 XI1.XI0.XI0.XI7<7>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<7>.MM_i_73 XI1.XI0.XI0.XI7<7>.NET_007
+ XI1.XI0.XI0.XI7<7>.NET_000 XI1.XI0.XI0.XI7<7>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<7>.MM_i_79 VDD! XI1.XI0.XI0.XI7<7>.NET_005
+ XI1.XI0.XI0.XI7<7>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<7>.MM_i_85 VDD! XI1.XI0.XI0.XI7<7>.NET_003
+ XI1.XI0.XI0.XI7<7>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<7>.MM_i_92 XI1.XI0.M_DATA<7> XI1.XI0.XI0.XI7<7>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<7>.MM_i_48 XI1.XI0.XI0.XI7<7>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<6>.MM_i_7 VSS! XI1.XI0.XI0.XI7<6>.NET_000
+ XI1.XI0.XI0.XI7<6>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<6>.MM_i_13 XI1.XI0.XI0.XI7<6>.NET_002 WR_DATA<6> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<6>.MM_i_18 XI1.XI0.XI0.XI7<6>.NET_003
+ XI1.XI0.XI0.XI7<6>.NET_000 XI1.XI0.XI0.XI7<6>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<6>.MM_i_24 XI1.XI0.XI0.XI7<6>.NET_004
+ XI1.XI0.XI0.XI7<6>.NET_001 XI1.XI0.XI0.XI7<6>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<6>.MM_i_29 VSS! XI1.XI0.XI0.XI7<6>.NET_005
+ XI1.XI0.XI0.XI7<6>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<6>.MM_i_35 VSS! XI1.XI0.XI0.XI7<6>.NET_003
+ XI1.XI0.XI0.XI7<6>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<6>.MM_i_42 XI1.XI0.M_DATA<6> XI1.XI0.XI0.XI7<6>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<6>.MM_i_0 XI1.XI0.XI0.XI7<6>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<6>.MM_i_55 VDD! XI1.XI0.XI0.XI7<6>.NET_000
+ XI1.XI0.XI0.XI7<6>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<6>.MM_i_62 XI1.XI0.XI0.XI7<6>.NET_006 WR_DATA<6> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<6>.MM_i_67 XI1.XI0.XI0.XI7<6>.NET_003
+ XI1.XI0.XI0.XI7<6>.NET_001 XI1.XI0.XI0.XI7<6>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<6>.MM_i_73 XI1.XI0.XI0.XI7<6>.NET_007
+ XI1.XI0.XI0.XI7<6>.NET_000 XI1.XI0.XI0.XI7<6>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<6>.MM_i_79 VDD! XI1.XI0.XI0.XI7<6>.NET_005
+ XI1.XI0.XI0.XI7<6>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<6>.MM_i_85 VDD! XI1.XI0.XI0.XI7<6>.NET_003
+ XI1.XI0.XI0.XI7<6>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<6>.MM_i_92 XI1.XI0.M_DATA<6> XI1.XI0.XI0.XI7<6>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<6>.MM_i_48 XI1.XI0.XI0.XI7<6>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<5>.MM_i_7 VSS! XI1.XI0.XI0.XI7<5>.NET_000
+ XI1.XI0.XI0.XI7<5>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<5>.MM_i_13 XI1.XI0.XI0.XI7<5>.NET_002 WR_DATA<5> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<5>.MM_i_18 XI1.XI0.XI0.XI7<5>.NET_003
+ XI1.XI0.XI0.XI7<5>.NET_000 XI1.XI0.XI0.XI7<5>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<5>.MM_i_24 XI1.XI0.XI0.XI7<5>.NET_004
+ XI1.XI0.XI0.XI7<5>.NET_001 XI1.XI0.XI0.XI7<5>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<5>.MM_i_29 VSS! XI1.XI0.XI0.XI7<5>.NET_005
+ XI1.XI0.XI0.XI7<5>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<5>.MM_i_35 VSS! XI1.XI0.XI0.XI7<5>.NET_003
+ XI1.XI0.XI0.XI7<5>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<5>.MM_i_42 XI1.XI0.M_DATA<5> XI1.XI0.XI0.XI7<5>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<5>.MM_i_0 XI1.XI0.XI0.XI7<5>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<5>.MM_i_55 VDD! XI1.XI0.XI0.XI7<5>.NET_000
+ XI1.XI0.XI0.XI7<5>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<5>.MM_i_62 XI1.XI0.XI0.XI7<5>.NET_006 WR_DATA<5> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<5>.MM_i_67 XI1.XI0.XI0.XI7<5>.NET_003
+ XI1.XI0.XI0.XI7<5>.NET_001 XI1.XI0.XI0.XI7<5>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<5>.MM_i_73 XI1.XI0.XI0.XI7<5>.NET_007
+ XI1.XI0.XI0.XI7<5>.NET_000 XI1.XI0.XI0.XI7<5>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<5>.MM_i_79 VDD! XI1.XI0.XI0.XI7<5>.NET_005
+ XI1.XI0.XI0.XI7<5>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<5>.MM_i_85 VDD! XI1.XI0.XI0.XI7<5>.NET_003
+ XI1.XI0.XI0.XI7<5>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<5>.MM_i_92 XI1.XI0.M_DATA<5> XI1.XI0.XI0.XI7<5>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<5>.MM_i_48 XI1.XI0.XI0.XI7<5>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<4>.MM_i_7 VSS! XI1.XI0.XI0.XI7<4>.NET_000
+ XI1.XI0.XI0.XI7<4>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<4>.MM_i_13 XI1.XI0.XI0.XI7<4>.NET_002 WR_DATA<4> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<4>.MM_i_18 XI1.XI0.XI0.XI7<4>.NET_003
+ XI1.XI0.XI0.XI7<4>.NET_000 XI1.XI0.XI0.XI7<4>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<4>.MM_i_24 XI1.XI0.XI0.XI7<4>.NET_004
+ XI1.XI0.XI0.XI7<4>.NET_001 XI1.XI0.XI0.XI7<4>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<4>.MM_i_29 VSS! XI1.XI0.XI0.XI7<4>.NET_005
+ XI1.XI0.XI0.XI7<4>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<4>.MM_i_35 VSS! XI1.XI0.XI0.XI7<4>.NET_003
+ XI1.XI0.XI0.XI7<4>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<4>.MM_i_42 XI1.XI0.M_DATA<4> XI1.XI0.XI0.XI7<4>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<4>.MM_i_0 XI1.XI0.XI0.XI7<4>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<4>.MM_i_55 VDD! XI1.XI0.XI0.XI7<4>.NET_000
+ XI1.XI0.XI0.XI7<4>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<4>.MM_i_62 XI1.XI0.XI0.XI7<4>.NET_006 WR_DATA<4> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<4>.MM_i_67 XI1.XI0.XI0.XI7<4>.NET_003
+ XI1.XI0.XI0.XI7<4>.NET_001 XI1.XI0.XI0.XI7<4>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<4>.MM_i_73 XI1.XI0.XI0.XI7<4>.NET_007
+ XI1.XI0.XI0.XI7<4>.NET_000 XI1.XI0.XI0.XI7<4>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<4>.MM_i_79 VDD! XI1.XI0.XI0.XI7<4>.NET_005
+ XI1.XI0.XI0.XI7<4>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<4>.MM_i_85 VDD! XI1.XI0.XI0.XI7<4>.NET_003
+ XI1.XI0.XI0.XI7<4>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<4>.MM_i_92 XI1.XI0.M_DATA<4> XI1.XI0.XI0.XI7<4>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<4>.MM_i_48 XI1.XI0.XI0.XI7<4>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<11>.MM_i_7 VSS! XI1.XI0.XI0.XI7<11>.NET_000
+ XI1.XI0.XI0.XI7<11>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<11>.MM_i_13 XI1.XI0.XI0.XI7<11>.NET_002 WR_DATA<11> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<11>.MM_i_18 XI1.XI0.XI0.XI7<11>.NET_003
+ XI1.XI0.XI0.XI7<11>.NET_000 XI1.XI0.XI0.XI7<11>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<11>.MM_i_24 XI1.XI0.XI0.XI7<11>.NET_004
+ XI1.XI0.XI0.XI7<11>.NET_001 XI1.XI0.XI0.XI7<11>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<11>.MM_i_29 VSS! XI1.XI0.XI0.XI7<11>.NET_005
+ XI1.XI0.XI0.XI7<11>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<11>.MM_i_35 VSS! XI1.XI0.XI0.XI7<11>.NET_003
+ XI1.XI0.XI0.XI7<11>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<11>.MM_i_42 XI1.XI0.M_DATA<11> XI1.XI0.XI0.XI7<11>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<11>.MM_i_0 XI1.XI0.XI0.XI7<11>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<11>.MM_i_55 VDD! XI1.XI0.XI0.XI7<11>.NET_000
+ XI1.XI0.XI0.XI7<11>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<11>.MM_i_62 XI1.XI0.XI0.XI7<11>.NET_006 WR_DATA<11> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<11>.MM_i_67 XI1.XI0.XI0.XI7<11>.NET_003
+ XI1.XI0.XI0.XI7<11>.NET_001 XI1.XI0.XI0.XI7<11>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<11>.MM_i_73 XI1.XI0.XI0.XI7<11>.NET_007
+ XI1.XI0.XI0.XI7<11>.NET_000 XI1.XI0.XI0.XI7<11>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<11>.MM_i_79 VDD! XI1.XI0.XI0.XI7<11>.NET_005
+ XI1.XI0.XI0.XI7<11>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<11>.MM_i_85 VDD! XI1.XI0.XI0.XI7<11>.NET_003
+ XI1.XI0.XI0.XI7<11>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<11>.MM_i_92 XI1.XI0.M_DATA<11> XI1.XI0.XI0.XI7<11>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<11>.MM_i_48 XI1.XI0.XI0.XI7<11>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<10>.MM_i_7 VSS! XI1.XI0.XI0.XI7<10>.NET_000
+ XI1.XI0.XI0.XI7<10>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<10>.MM_i_13 XI1.XI0.XI0.XI7<10>.NET_002 WR_DATA<10> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<10>.MM_i_18 XI1.XI0.XI0.XI7<10>.NET_003
+ XI1.XI0.XI0.XI7<10>.NET_000 XI1.XI0.XI0.XI7<10>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<10>.MM_i_24 XI1.XI0.XI0.XI7<10>.NET_004
+ XI1.XI0.XI0.XI7<10>.NET_001 XI1.XI0.XI0.XI7<10>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<10>.MM_i_29 VSS! XI1.XI0.XI0.XI7<10>.NET_005
+ XI1.XI0.XI0.XI7<10>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<10>.MM_i_35 VSS! XI1.XI0.XI0.XI7<10>.NET_003
+ XI1.XI0.XI0.XI7<10>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<10>.MM_i_42 XI1.XI0.M_DATA<10> XI1.XI0.XI0.XI7<10>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<10>.MM_i_0 XI1.XI0.XI0.XI7<10>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<10>.MM_i_55 VDD! XI1.XI0.XI0.XI7<10>.NET_000
+ XI1.XI0.XI0.XI7<10>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<10>.MM_i_62 XI1.XI0.XI0.XI7<10>.NET_006 WR_DATA<10> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<10>.MM_i_67 XI1.XI0.XI0.XI7<10>.NET_003
+ XI1.XI0.XI0.XI7<10>.NET_001 XI1.XI0.XI0.XI7<10>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<10>.MM_i_73 XI1.XI0.XI0.XI7<10>.NET_007
+ XI1.XI0.XI0.XI7<10>.NET_000 XI1.XI0.XI0.XI7<10>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<10>.MM_i_79 VDD! XI1.XI0.XI0.XI7<10>.NET_005
+ XI1.XI0.XI0.XI7<10>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<10>.MM_i_85 VDD! XI1.XI0.XI0.XI7<10>.NET_003
+ XI1.XI0.XI0.XI7<10>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<10>.MM_i_92 XI1.XI0.M_DATA<10> XI1.XI0.XI0.XI7<10>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<10>.MM_i_48 XI1.XI0.XI0.XI7<10>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<9>.MM_i_7 VSS! XI1.XI0.XI0.XI7<9>.NET_000
+ XI1.XI0.XI0.XI7<9>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<9>.MM_i_13 XI1.XI0.XI0.XI7<9>.NET_002 WR_DATA<9> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<9>.MM_i_18 XI1.XI0.XI0.XI7<9>.NET_003
+ XI1.XI0.XI0.XI7<9>.NET_000 XI1.XI0.XI0.XI7<9>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<9>.MM_i_24 XI1.XI0.XI0.XI7<9>.NET_004
+ XI1.XI0.XI0.XI7<9>.NET_001 XI1.XI0.XI0.XI7<9>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<9>.MM_i_29 VSS! XI1.XI0.XI0.XI7<9>.NET_005
+ XI1.XI0.XI0.XI7<9>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<9>.MM_i_35 VSS! XI1.XI0.XI0.XI7<9>.NET_003
+ XI1.XI0.XI0.XI7<9>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<9>.MM_i_42 XI1.XI0.M_DATA<9> XI1.XI0.XI0.XI7<9>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<9>.MM_i_0 XI1.XI0.XI0.XI7<9>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<9>.MM_i_55 VDD! XI1.XI0.XI0.XI7<9>.NET_000
+ XI1.XI0.XI0.XI7<9>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<9>.MM_i_62 XI1.XI0.XI0.XI7<9>.NET_006 WR_DATA<9> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<9>.MM_i_67 XI1.XI0.XI0.XI7<9>.NET_003
+ XI1.XI0.XI0.XI7<9>.NET_001 XI1.XI0.XI0.XI7<9>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<9>.MM_i_73 XI1.XI0.XI0.XI7<9>.NET_007
+ XI1.XI0.XI0.XI7<9>.NET_000 XI1.XI0.XI0.XI7<9>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<9>.MM_i_79 VDD! XI1.XI0.XI0.XI7<9>.NET_005
+ XI1.XI0.XI0.XI7<9>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<9>.MM_i_85 VDD! XI1.XI0.XI0.XI7<9>.NET_003
+ XI1.XI0.XI0.XI7<9>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<9>.MM_i_92 XI1.XI0.M_DATA<9> XI1.XI0.XI0.XI7<9>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<9>.MM_i_48 XI1.XI0.XI0.XI7<9>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<8>.MM_i_7 VSS! XI1.XI0.XI0.XI7<8>.NET_000
+ XI1.XI0.XI0.XI7<8>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<8>.MM_i_13 XI1.XI0.XI0.XI7<8>.NET_002 WR_DATA<8> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<8>.MM_i_18 XI1.XI0.XI0.XI7<8>.NET_003
+ XI1.XI0.XI0.XI7<8>.NET_000 XI1.XI0.XI0.XI7<8>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<8>.MM_i_24 XI1.XI0.XI0.XI7<8>.NET_004
+ XI1.XI0.XI0.XI7<8>.NET_001 XI1.XI0.XI0.XI7<8>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<8>.MM_i_29 VSS! XI1.XI0.XI0.XI7<8>.NET_005
+ XI1.XI0.XI0.XI7<8>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<8>.MM_i_35 VSS! XI1.XI0.XI0.XI7<8>.NET_003
+ XI1.XI0.XI0.XI7<8>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<8>.MM_i_42 XI1.XI0.M_DATA<8> XI1.XI0.XI0.XI7<8>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<8>.MM_i_0 XI1.XI0.XI0.XI7<8>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<8>.MM_i_55 VDD! XI1.XI0.XI0.XI7<8>.NET_000
+ XI1.XI0.XI0.XI7<8>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<8>.MM_i_62 XI1.XI0.XI0.XI7<8>.NET_006 WR_DATA<8> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<8>.MM_i_67 XI1.XI0.XI0.XI7<8>.NET_003
+ XI1.XI0.XI0.XI7<8>.NET_001 XI1.XI0.XI0.XI7<8>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<8>.MM_i_73 XI1.XI0.XI0.XI7<8>.NET_007
+ XI1.XI0.XI0.XI7<8>.NET_000 XI1.XI0.XI0.XI7<8>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<8>.MM_i_79 VDD! XI1.XI0.XI0.XI7<8>.NET_005
+ XI1.XI0.XI0.XI7<8>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<8>.MM_i_85 VDD! XI1.XI0.XI0.XI7<8>.NET_003
+ XI1.XI0.XI0.XI7<8>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<8>.MM_i_92 XI1.XI0.M_DATA<8> XI1.XI0.XI0.XI7<8>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<8>.MM_i_48 XI1.XI0.XI0.XI7<8>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<15>.MM_i_7 VSS! XI1.XI0.XI0.XI7<15>.NET_000
+ XI1.XI0.XI0.XI7<15>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<15>.MM_i_13 XI1.XI0.XI0.XI7<15>.NET_002 WR_DATA<15> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<15>.MM_i_18 XI1.XI0.XI0.XI7<15>.NET_003
+ XI1.XI0.XI0.XI7<15>.NET_000 XI1.XI0.XI0.XI7<15>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<15>.MM_i_24 XI1.XI0.XI0.XI7<15>.NET_004
+ XI1.XI0.XI0.XI7<15>.NET_001 XI1.XI0.XI0.XI7<15>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<15>.MM_i_29 VSS! XI1.XI0.XI0.XI7<15>.NET_005
+ XI1.XI0.XI0.XI7<15>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<15>.MM_i_35 VSS! XI1.XI0.XI0.XI7<15>.NET_003
+ XI1.XI0.XI0.XI7<15>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<15>.MM_i_42 XI1.XI0.M_DATA<15> XI1.XI0.XI0.XI7<15>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<15>.MM_i_0 XI1.XI0.XI0.XI7<15>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<15>.MM_i_55 VDD! XI1.XI0.XI0.XI7<15>.NET_000
+ XI1.XI0.XI0.XI7<15>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<15>.MM_i_62 XI1.XI0.XI0.XI7<15>.NET_006 WR_DATA<15> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<15>.MM_i_67 XI1.XI0.XI0.XI7<15>.NET_003
+ XI1.XI0.XI0.XI7<15>.NET_001 XI1.XI0.XI0.XI7<15>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<15>.MM_i_73 XI1.XI0.XI0.XI7<15>.NET_007
+ XI1.XI0.XI0.XI7<15>.NET_000 XI1.XI0.XI0.XI7<15>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<15>.MM_i_79 VDD! XI1.XI0.XI0.XI7<15>.NET_005
+ XI1.XI0.XI0.XI7<15>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<15>.MM_i_85 VDD! XI1.XI0.XI0.XI7<15>.NET_003
+ XI1.XI0.XI0.XI7<15>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<15>.MM_i_92 XI1.XI0.M_DATA<15> XI1.XI0.XI0.XI7<15>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<15>.MM_i_48 XI1.XI0.XI0.XI7<15>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<14>.MM_i_7 VSS! XI1.XI0.XI0.XI7<14>.NET_000
+ XI1.XI0.XI0.XI7<14>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<14>.MM_i_13 XI1.XI0.XI0.XI7<14>.NET_002 WR_DATA<14> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<14>.MM_i_18 XI1.XI0.XI0.XI7<14>.NET_003
+ XI1.XI0.XI0.XI7<14>.NET_000 XI1.XI0.XI0.XI7<14>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<14>.MM_i_24 XI1.XI0.XI0.XI7<14>.NET_004
+ XI1.XI0.XI0.XI7<14>.NET_001 XI1.XI0.XI0.XI7<14>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<14>.MM_i_29 VSS! XI1.XI0.XI0.XI7<14>.NET_005
+ XI1.XI0.XI0.XI7<14>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<14>.MM_i_35 VSS! XI1.XI0.XI0.XI7<14>.NET_003
+ XI1.XI0.XI0.XI7<14>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<14>.MM_i_42 XI1.XI0.M_DATA<14> XI1.XI0.XI0.XI7<14>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<14>.MM_i_0 XI1.XI0.XI0.XI7<14>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<14>.MM_i_55 VDD! XI1.XI0.XI0.XI7<14>.NET_000
+ XI1.XI0.XI0.XI7<14>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<14>.MM_i_62 XI1.XI0.XI0.XI7<14>.NET_006 WR_DATA<14> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<14>.MM_i_67 XI1.XI0.XI0.XI7<14>.NET_003
+ XI1.XI0.XI0.XI7<14>.NET_001 XI1.XI0.XI0.XI7<14>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<14>.MM_i_73 XI1.XI0.XI0.XI7<14>.NET_007
+ XI1.XI0.XI0.XI7<14>.NET_000 XI1.XI0.XI0.XI7<14>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<14>.MM_i_79 VDD! XI1.XI0.XI0.XI7<14>.NET_005
+ XI1.XI0.XI0.XI7<14>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<14>.MM_i_85 VDD! XI1.XI0.XI0.XI7<14>.NET_003
+ XI1.XI0.XI0.XI7<14>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<14>.MM_i_92 XI1.XI0.M_DATA<14> XI1.XI0.XI0.XI7<14>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<14>.MM_i_48 XI1.XI0.XI0.XI7<14>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<13>.MM_i_7 VSS! XI1.XI0.XI0.XI7<13>.NET_000
+ XI1.XI0.XI0.XI7<13>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<13>.MM_i_13 XI1.XI0.XI0.XI7<13>.NET_002 WR_DATA<13> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<13>.MM_i_18 XI1.XI0.XI0.XI7<13>.NET_003
+ XI1.XI0.XI0.XI7<13>.NET_000 XI1.XI0.XI0.XI7<13>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<13>.MM_i_24 XI1.XI0.XI0.XI7<13>.NET_004
+ XI1.XI0.XI0.XI7<13>.NET_001 XI1.XI0.XI0.XI7<13>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<13>.MM_i_29 VSS! XI1.XI0.XI0.XI7<13>.NET_005
+ XI1.XI0.XI0.XI7<13>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<13>.MM_i_35 VSS! XI1.XI0.XI0.XI7<13>.NET_003
+ XI1.XI0.XI0.XI7<13>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<13>.MM_i_42 XI1.XI0.M_DATA<13> XI1.XI0.XI0.XI7<13>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<13>.MM_i_0 XI1.XI0.XI0.XI7<13>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<13>.MM_i_55 VDD! XI1.XI0.XI0.XI7<13>.NET_000
+ XI1.XI0.XI0.XI7<13>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<13>.MM_i_62 XI1.XI0.XI0.XI7<13>.NET_006 WR_DATA<13> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<13>.MM_i_67 XI1.XI0.XI0.XI7<13>.NET_003
+ XI1.XI0.XI0.XI7<13>.NET_001 XI1.XI0.XI0.XI7<13>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<13>.MM_i_73 XI1.XI0.XI0.XI7<13>.NET_007
+ XI1.XI0.XI0.XI7<13>.NET_000 XI1.XI0.XI0.XI7<13>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<13>.MM_i_79 VDD! XI1.XI0.XI0.XI7<13>.NET_005
+ XI1.XI0.XI0.XI7<13>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<13>.MM_i_85 VDD! XI1.XI0.XI0.XI7<13>.NET_003
+ XI1.XI0.XI0.XI7<13>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<13>.MM_i_92 XI1.XI0.M_DATA<13> XI1.XI0.XI0.XI7<13>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<13>.MM_i_48 XI1.XI0.XI0.XI7<13>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI0.XI7<12>.MM_i_7 VSS! XI1.XI0.XI0.XI7<12>.NET_000
+ XI1.XI0.XI0.XI7<12>.NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI1.XI0.XI0.XI7<12>.MM_i_13 XI1.XI0.XI0.XI7<12>.NET_002 WR_DATA<12> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<12>.MM_i_18 XI1.XI0.XI0.XI7<12>.NET_003
+ XI1.XI0.XI0.XI7<12>.NET_000 XI1.XI0.XI0.XI7<12>.NET_002 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.145e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI1.XI0.XI0.XI7<12>.MM_i_24 XI1.XI0.XI0.XI7<12>.NET_004
+ XI1.XI0.XI0.XI7<12>.NET_001 XI1.XI0.XI0.XI7<12>.NET_003 VSS! NMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.145e-14 PD=4.6e-07 PS=7e-07
mXI1.XI0.XI0.XI7<12>.MM_i_29 VSS! XI1.XI0.XI0.XI7<12>.NET_005
+ XI1.XI0.XI0.XI7<12>.NET_004 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<12>.MM_i_35 VSS! XI1.XI0.XI0.XI7<12>.NET_003
+ XI1.XI0.XI0.XI7<12>.NET_005 VSS! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<12>.MM_i_42 XI1.XI0.M_DATA<12> XI1.XI0.XI0.XI7<12>.NET_003 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI1.XI0.XI0.XI7<12>.MM_i_0 XI1.XI0.XI0.XI7<12>.NET_000 XI1.XI0.CLK_N VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=4.375e-14 PD=6.3e-07 PS=1.11e-06
mXI1.XI0.XI0.XI7<12>.MM_i_55 VDD! XI1.XI0.XI0.XI7<12>.NET_000
+ XI1.XI0.XI0.XI7<12>.NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI1.XI0.XI0.XI7<12>.MM_i_62 XI1.XI0.XI0.XI7<12>.NET_006 WR_DATA<12> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<12>.MM_i_67 XI1.XI0.XI0.XI7<12>.NET_003
+ XI1.XI0.XI0.XI7<12>.NET_001 XI1.XI0.XI0.XI7<12>.NET_006 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=2.855e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<12>.MM_i_73 XI1.XI0.XI0.XI7<12>.NET_007
+ XI1.XI0.XI0.XI7<12>.NET_000 XI1.XI0.XI0.XI7<12>.NET_003 VDD! PMOS_VTL L=5e-08
+ W=9e-08 AD=1.26e-14 AS=2.855e-14 PD=4.6e-07 PS=9.1e-07
mXI1.XI0.XI0.XI7<12>.MM_i_79 VDD! XI1.XI0.XI0.XI7<12>.NET_005
+ XI1.XI0.XI0.XI7<12>.NET_007 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=1.26e-14 PD=4.6e-07 PS=4.6e-07
mXI1.XI0.XI0.XI7<12>.MM_i_85 VDD! XI1.XI0.XI0.XI7<12>.NET_003
+ XI1.XI0.XI0.XI7<12>.NET_005 VDD! PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14
+ AS=9.45e-15 PD=4.6e-07 PS=3.9e-07
mXI1.XI0.XI0.XI7<12>.MM_i_92 XI1.XI0.M_DATA<12> XI1.XI0.XI0.XI7<12>.NET_003 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI1.XI0.XI0.XI7<12>.MM_i_48 XI1.XI0.XI0.XI7<12>.NET_000 XI1.XI0.CLK_N VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06
mXI1.XI0.XI21<1>.MM_i_2 VSS! CLK XI1.XI0.XI21<1>.Z_NEG VSS! NMOS_VTL L=5e-08
+ W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI21<1>.MM_i_0_0 VSS! XI1.XI0.XI21<1>.Z_NEG XI1.XI0.CK VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07
mXI1.XI0.XI21<1>.MM_i_0_1 VSS! XI1.XI0.XI21<1>.Z_NEG XI1.XI0.CK VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07
mXI1.XI0.XI21<1>.MM_i_3 VDD! CLK XI1.XI0.XI21<1>.Z_NEG VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI21<1>.MM_i_1_0 VDD! XI1.XI0.XI21<1>.Z_NEG XI1.XI0.CK VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI21<1>.MM_i_1_1 VDD! XI1.XI0.XI21<1>.Z_NEG XI1.XI0.CK VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI21<0>.MM_i_2 VSS! CLK XI1.XI0.XI21<0>.Z_NEG VSS! NMOS_VTL L=5e-08
+ W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI21<0>.MM_i_0_0 VSS! XI1.XI0.XI21<0>.Z_NEG XI1.XI0.CK VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07
mXI1.XI0.XI21<0>.MM_i_0_1 VSS! XI1.XI0.XI21<0>.Z_NEG XI1.XI0.CK VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07
mXI1.XI0.XI21<0>.MM_i_3 VDD! CLK XI1.XI0.XI21<0>.Z_NEG VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI21<0>.MM_i_1_0 VDD! XI1.XI0.XI21<0>.Z_NEG XI1.XI0.CK VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI21<0>.MM_i_1_1 VDD! XI1.XI0.XI21<0>.Z_NEG XI1.XI0.CK VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI1.XI0.XI20.MM_i_2 VSS! XI1.XI0.CLK_PREBUFF XI1.XI0.XI20.Z_NEG VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07
mXI1.XI0.XI20.MM_i_0_0 VSS! XI1.XI0.XI20.Z_NEG XI1.XI0.CLK_N VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07
mXI1.XI0.XI20.MM_i_0_1 VSS! XI1.XI0.XI20.Z_NEG XI1.XI0.CLK_N VSS! NMOS_VTL
+ L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07
mXI1.XI0.XI20.MM_i_3 VDD! XI1.XI0.CLK_PREBUFF XI1.XI0.XI20.Z_NEG VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI1.XI0.XI20.MM_i_1_0 VDD! XI1.XI0.XI20.Z_NEG XI1.XI0.CLK_N VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI1.XI0.XI20.MM_i_1_1 VDD! XI1.XI0.XI20.Z_NEG XI1.XI0.CLK_N VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
c_2217 VDD! 0 120.767f
c_4434 VSS! 0 116.598f
c_4444 WR_DATA<4> 0 0.0408626f
c_4454 WR_DATA<6> 0 0.0408626f
c_4464 WR_DATA<1> 0 0.0408626f
c_4474 WR_DATA<2> 0 0.0408626f
c_4484 WR_DATA<11> 0 0.0408626f
c_4494 WR_DATA<12> 0 0.0411361f
c_4504 WR_DATA<15> 0 0.0410413f
c_4514 WR_DATA<0> 0 0.0409312f
c_4524 WR_DATA<13> 0 0.0408491f
c_4534 WR_DATA<14> 0 0.0408626f
c_4544 WR_DATA<8> 0 0.0409312f
c_4554 WR_DATA<9> 0 0.0408626f
c_4564 WR_DATA<3> 0 0.0408626f
c_4574 WR_DATA<10> 0 0.0408626f
c_4584 WR_DATA<5> 0 0.0408626f
c_4594 WR_DATA<7> 0 0.0409312f
c_4918 REG_DATA_11<9> 0 1.22983f
c_5016 RD_DATA_0<8> 0 0.609292f
c_5092 RD_DATA_0<3> 0 0.598651f
c_5209 RD_DATA_0<12> 0 0.601737f
c_5289 RD_DATA_0<4> 0 0.612548f
c_5379 RD_DATA_0<6> 0 0.610717f
c_5508 RD_DATA_0<14> 0 0.519789f
c_5611 RD_DATA_0<9> 0 0.592099f
c_5689 RD_DATA_0<0> 0 0.618411f
c_5797 RD_DATA_0<10> 0 0.608483f
c_5867 RD_DATA_0<2> 0 0.653963f
c_5981 RD_DATA_0<11> 0 0.590637f
c_6113 RD_DATA_0<15> 0 0.490872f
c_6207 RD_DATA_0<7> 0 0.588356f
c_6335 RD_DATA_0<13> 0 0.582146f
c_6420 RD_DATA_0<5> 0 0.593781f
c_6487 RD_DATA_0<1> 0 0.599491f
c_6563 REG_DATA_0<0> 0 3.62623f
c_6639 REG_DATA_1<0> 0 1.0436f
c_6715 REG_DATA_2<0> 0 1.64217f
c_6791 REG_DATA_3<0> 0 1.73139f
c_6867 REG_DATA_4<0> 0 1.8742f
c_6943 REG_DATA_5<0> 0 1.9455f
c_7020 REG_DATA_6<0> 0 1.86013f
c_7097 REG_DATA_7<0> 0 1.77272f
c_7198 REG_DATA_8<0> 0 1.42434f
c_7299 REG_DATA_9<0> 0 1.41631f
c_7448 REG_DATA_10<0> 0 1.6055f
c_7597 REG_DATA_11<0> 0 1.19582f
c_7770 REG_DATA_12<0> 0 1.73017f
c_7957 REG_DATA_0<1> 0 1.66633f
c_8146 REG_DATA_1<1> 0 1.66612f
c_8313 REG_DATA_2<1> 0 1.77856f
c_8478 REG_DATA_3<1> 0 1.57539f
c_8643 REG_DATA_4<1> 0 1.43982f
c_8806 REG_DATA_5<1> 0 1.6838f
c_8971 REG_DATA_6<1> 0 1.59782f
c_9158 REG_DATA_7<1> 0 1.60026f
c_9345 REG_DATA_8<1> 0 1.20856f
c_9508 REG_DATA_9<1> 0 1.53846f
c_9671 REG_DATA_10<1> 0 1.65976f
c_9836 REG_DATA_11<1> 0 1.44516f
c_9948 REG_DATA_12<1> 0 1.36729f
c_10113 REG_DATA_0<2> 0 1.80067f
c_10278 REG_DATA_1<2> 0 1.97486f
c_10469 REG_DATA_2<2> 0 1.87514f
c_10658 REG_DATA_3<2> 0 1.94591f
c_10847 REG_DATA_4<2> 0 2.09173f
c_11021 REG_DATA_5<2> 0 1.90752f
c_11195 REG_DATA_6<2> 0 1.90258f
c_11369 REG_DATA_7<2> 0 1.84686f
c_11545 REG_DATA_8<2> 0 2.21902f
c_11723 REG_DATA_9<2> 0 2.25676f
c_11925 REG_DATA_10<2> 0 2.22083f
c_12127 REG_DATA_11<2> 0 2.24387f
c_12304 REG_DATA_12<2> 0 1.97922f
c_12484 REG_DATA_0<3> 0 2.11736f
c_12680 REG_DATA_1<3> 0 1.85975f
c_12834 REG_DATA_2<3> 0 1.58998f
c_13036 REG_DATA_3<3> 0 2.10534f
c_13240 REG_DATA_4<3> 0 2.26143f
c_13470 REG_DATA_5<3> 0 2.36641f
c_13701 REG_DATA_6<3> 0 2.08525f
c_13933 REG_DATA_7<3> 0 2.03275f
c_14152 REG_DATA_8<3> 0 2.06143f
c_14363 REG_DATA_9<3> 0 1.79091f
c_14582 REG_DATA_10<3> 0 1.6868f
c_14801 REG_DATA_11<3> 0 1.83712f
c_15047 REG_DATA_12<3> 0 1.84349f
c_15351 REG_DATA_0<4> 0 2.1204f
c_15656 REG_DATA_1<4> 0 1.64671f
c_15936 REG_DATA_2<4> 0 1.55707f
c_16216 REG_DATA_3<4> 0 1.90758f
c_16499 REG_DATA_4<4> 0 1.47116f
c_16731 REG_DATA_5<4> 0 1.24556f
c_16954 REG_DATA_6<4> 0 1.27865f
c_17224 REG_DATA_7<4> 0 1.56751f
c_17522 REG_DATA_8<4> 0 1.6971f
c_17821 REG_DATA_9<4> 0 1.9941f
c_18120 REG_DATA_10<4> 0 1.5066f
c_18399 REG_DATA_11<4> 0 1.36783f
c_18665 REG_DATA_12<4> 0 1.19282f
c_18916 REG_DATA_0<5> 0 0.922496f
c_19178 REG_DATA_1<5> 0 1.48207f
c_19448 REG_DATA_2<5> 0 1.92198f
c_19735 REG_DATA_3<5> 0 1.93075f
c_20022 REG_DATA_4<5> 0 2.18569f
c_20284 REG_DATA_5<5> 0 1.70824f
c_20545 REG_DATA_6<5> 0 1.57214f
c_20753 REG_DATA_7<5> 0 1.14585f
c_20959 REG_DATA_8<5> 0 1.23743f
c_21230 REG_DATA_9<5> 0 1.5433f
c_21501 REG_DATA_10<5> 0 2.01145f
c_21798 REG_DATA_11<5> 0 1.82128f
c_22086 REG_DATA_12<5> 0 1.59599f
c_22367 REG_DATA_0<6> 0 1.39177f
c_22624 REG_DATA_1<6> 0 1.25786f
c_22880 REG_DATA_2<6> 0 1.23081f
c_23137 REG_DATA_3<6> 0 1.11949f
c_23408 REG_DATA_4<6> 0 1.45033f
c_23681 REG_DATA_5<6> 0 1.97452f
c_23975 REG_DATA_6<6> 0 1.74777f
c_24267 REG_DATA_7<6> 0 1.80032f
c_24485 REG_DATA_8<6> 0 1.32493f
c_24751 REG_DATA_9<6> 0 1.57325f
c_25020 REG_DATA_10<6> 0 1.3354f
c_25239 REG_DATA_11<6> 0 1.58485f
c_25522 REG_DATA_12<6> 0 1.54964f
c_25792 REG_DATA_0<7> 0 1.51807f
c_26093 REG_DATA_1<7> 0 1.75029f
c_26387 REG_DATA_2<7> 0 1.39972f
c_26683 REG_DATA_3<7> 0 1.52227f
c_26960 REG_DATA_4<7> 0 1.67598f
c_27235 REG_DATA_5<7> 0 1.35622f
c_27513 REG_DATA_6<7> 0 1.55463f
c_27803 REG_DATA_7<7> 0 1.68937f
c_28082 REG_DATA_8<7> 0 1.65046f
c_28334 REG_DATA_9<7> 0 1.66523f
c_28635 REG_DATA_10<7> 0 1.78692f
c_28911 REG_DATA_11<7> 0 1.58618f
c_29188 REG_DATA_12<7> 0 2.04839f
c_29455 REG_DATA_0<8> 0 1.49214f
c_29677 REG_DATA_1<8> 0 1.14912f
c_29963 REG_DATA_2<8> 0 1.5035f
c_30221 REG_DATA_3<8> 0 1.27876f
c_30479 REG_DATA_4<8> 0 1.90633f
c_30738 REG_DATA_5<8> 0 1.97857f
c_30996 REG_DATA_6<8> 0 1.71968f
c_31233 REG_DATA_7<8> 0 1.75786f
c_31471 REG_DATA_8<8> 0 1.53791f
c_31706 REG_DATA_9<8> 0 1.39322f
c_31955 REG_DATA_10<8> 0 1.70763f
c_32206 REG_DATA_11<8> 0 1.87359f
c_32478 REG_DATA_12<8> 0 1.84796f
c_32738 REG_DATA_0<9> 0 1.51529f
c_32985 REG_DATA_1<9> 0 1.64987f
c_33232 REG_DATA_2<9> 0 1.71047f
c_33479 REG_DATA_3<9> 0 1.65768f
c_33742 REG_DATA_4<9> 0 1.13126f
c_34046 REG_DATA_5<9> 0 1.23201f
c_34369 REG_DATA_6<9> 0 1.48515f
c_34716 REG_DATA_7<9> 0 1.72661f
c_35063 REG_DATA_8<9> 0 1.6446f
c_35410 REG_DATA_9<9> 0 1.9967f
c_35737 REG_DATA_10<9> 0 1.68361f
c_36015 REG_DATA_12<9> 0 0.782248f
c_36329 REG_DATA_0<10> 0 1.48969f
c_36654 REG_DATA_1<10> 0 1.61202f
c_37002 REG_DATA_2<10> 0 2.23691f
c_37350 REG_DATA_3<10> 0 1.78924f
c_37672 REG_DATA_4<10> 0 1.5486f
c_37992 REG_DATA_5<10> 0 1.5666f
c_38310 REG_DATA_6<10> 0 1.08506f
c_38583 REG_DATA_7<10> 0 1.09184f
c_38856 REG_DATA_8<10> 0 1.2952f
c_39129 REG_DATA_9<10> 0 1.40799f
c_39402 REG_DATA_10<10> 0 1.93686f
c_39673 REG_DATA_11<10> 0 1.63367f
c_39936 REG_DATA_12<10> 0 1.55511f
c_40139 REG_DATA_0<11> 0 1.33618f
c_40398 REG_DATA_1<11> 0 1.46794f
c_40658 REG_DATA_2<11> 0 1.36331f
c_40917 REG_DATA_3<11> 0 1.38363f
c_41176 REG_DATA_4<11> 0 0.782461f
c_41435 REG_DATA_5<11> 0 1.22037f
c_41694 REG_DATA_6<11> 0 1.31179f
c_41949 REG_DATA_7<11> 0 1.27244f
c_42209 REG_DATA_8<11> 0 1.54922f
c_42470 REG_DATA_9<11> 0 1.54917f
c_42731 REG_DATA_10<11> 0 1.61663f
c_42990 REG_DATA_11<11> 0 1.82694f
c_43249 REG_DATA_12<11> 0 1.46173f
c_43449 REG_DATA_0<12> 0 0.730892f
c_43700 REG_DATA_1<12> 0 0.719026f
c_43951 REG_DATA_2<12> 0 1.2432f
c_44202 REG_DATA_3<12> 0 1.66223f
c_44453 REG_DATA_4<12> 0 1.56077f
c_44704 REG_DATA_5<12> 0 1.5236f
c_44956 REG_DATA_6<12> 0 1.53039f
c_45204 REG_DATA_7<12> 0 1.31918f
c_45454 REG_DATA_8<12> 0 1.42834f
c_45705 REG_DATA_9<12> 0 1.30458f
c_45956 REG_DATA_10<12> 0 0.966471f
c_46207 REG_DATA_11<12> 0 1.02312f
c_46455 REG_DATA_12<12> 0 1.27893f
c_46685 REG_DATA_0<13> 0 1.37356f
c_46871 REG_DATA_1<13> 0 1.3588f
c_47106 REG_DATA_2<13> 0 1.64295f
c_47342 REG_DATA_3<13> 0 1.63112f
c_47578 REG_DATA_4<13> 0 1.93626f
c_47814 REG_DATA_5<13> 0 1.49304f
c_48050 REG_DATA_6<13> 0 1.34097f
c_48284 REG_DATA_7<13> 0 0.878821f
c_48491 REG_DATA_8<13> 0 0.502049f
c_48674 REG_DATA_9<13> 0 1.17557f
c_48842 REG_DATA_10<13> 0 1.33358f
c_49010 REG_DATA_11<13> 0 1.6513f
c_49178 REG_DATA_12<13> 0 1.68546f
c_49331 REG_DATA_0<14> 0 1.95461f
c_49484 REG_DATA_1<14> 0 1.95199f
c_49637 REG_DATA_2<14> 0 1.74721f
c_49790 REG_DATA_3<14> 0 1.5589f
c_49943 REG_DATA_4<14> 0 1.05575f
c_50095 REG_DATA_5<14> 0 0.631894f
c_50247 REG_DATA_6<14> 0 1.44778f
c_50399 REG_DATA_7<14> 0 1.56108f
c_50551 REG_DATA_8<14> 0 1.87246f
c_50703 REG_DATA_9<14> 0 1.95206f
c_50855 REG_DATA_10<14> 0 1.95206f
c_51007 REG_DATA_11<14> 0 1.93928f
c_51156 REG_DATA_12<14> 0 1.71227f
c_51286 REG_DATA_0<15> 0 1.46512f
c_51418 REG_DATA_1<15> 0 0.904388f
c_51550 REG_DATA_2<15> 0 0.463885f
c_51682 REG_DATA_3<15> 0 1.33462f
c_51814 REG_DATA_4<15> 0 1.47114f
c_51946 REG_DATA_5<15> 0 1.7984f
c_52078 REG_DATA_6<15> 0 1.81264f
c_52210 REG_DATA_7<15> 0 1.8041f
c_52342 REG_DATA_8<15> 0 1.83706f
c_52474 REG_DATA_9<15> 0 1.64257f
c_52606 REG_DATA_10<15> 0 1.46957f
c_52738 REG_DATA_11<15> 0 0.895701f
c_52870 REG_DATA_12<15> 0 0.46986f
c_52968 RD_DATA_1<8> 0 0.609292f
c_53044 RD_DATA_1<3> 0 0.598651f
c_53161 RD_DATA_1<12> 0 0.601737f
c_53241 RD_DATA_1<4> 0 0.612548f
c_53331 RD_DATA_1<6> 0 0.610717f
c_53460 RD_DATA_1<14> 0 0.519789f
c_53563 RD_DATA_1<9> 0 0.592099f
c_53641 RD_DATA_1<0> 0 0.618411f
c_53749 RD_DATA_1<10> 0 0.608483f
c_53819 RD_DATA_1<2> 0 0.653963f
c_53933 RD_DATA_1<11> 0 0.590637f
c_54065 RD_DATA_1<15> 0 0.490872f
c_54159 RD_DATA_1<7> 0 0.588356f
c_54287 RD_DATA_1<13> 0 0.582146f
c_54372 RD_DATA_1<5> 0 0.593781f
c_54439 RD_DATA_1<1> 0 0.599491f
c_54473 CLK 0 0.767274f
c_54488 RD_ADDR_0<2> 0 0.758629f
c_54508 RD_ADDR_0<0> 0 0.893563f
c_54524 RD_ADDR_0<3> 0 1.03565f
c_54542 RD_ADDR_0<1> 0 0.672294f
c_54557 RD_ADDR_1<2> 0 0.745998f
c_54577 RD_ADDR_1<0> 0 0.790288f
c_54593 RD_ADDR_1<3> 0 0.928235f
c_54611 RD_ADDR_1<1> 0 0.665903f
c_54627 WR_ADDR<2> 0 0.758188f
c_54648 WR_ADDR<0> 0 0.892361f
c_54664 WR_EN 0 0.241236f
c_54681 WR_ADDR<3> 0 1.03449f
c_54700 WR_ADDR<1> 0 0.671853f
c_54969 XI0.NET1<0> 0 4.4071f
c_55238 XI0.NET1<1> 0 4.40746f
c_55508 XI0.NET1<2> 0 4.43707f
c_55779 XI0.NET1<3> 0 4.47328f
c_56052 XI0.NET1<4> 0 4.45238f
c_56325 XI0.NET1<5> 0 4.47808f
c_56600 XI0.NET1<6> 0 4.51347f
c_56874 XI0.NET1<7> 0 4.51618f
c_57151 XI0.NET1<8> 0 4.5833f
c_57429 XI0.NET1<9> 0 4.53587f
c_57704 XI0.NET1<10> 0 4.49353f
c_57978 XI0.NET1<11> 0 4.66969f
c_58235 XI0.NET1<12> 0 4.71897f
c_58243 XI0.XI0.NET_11XX 0 0.15093f
c_58274 XI0.XI0.NET_XX00 0 1.10722f
c_58296 XI0.XI0.NET_XX11 0 0.707171f
c_58313 XI0.XI0.NET_10XX 0 0.637717f
c_58329 XI0.XI0.ADDR_BAR<2> 0 0.648803f
c_58346 XI0.XI0.ADDR_BAR<0> 0 0.708334f
c_58370 XI0.XI0.NET_XX10 0 0.981965f
c_58388 XI0.XI0.NET_01XX 0 0.614487f
c_58403 XI0.XI0.ADDR_BAR<1> 0 0.524568f
c_58424 XI0.XI0.NET_XX01 0 0.972175f
c_58441 XI0.XI0.NET_00XX 0 0.630231f
c_58458 XI0.XI0.ADDR_BAR<3> 0 0.394208f
c_58465 XI0.XI0.XI11.ZN_NEG 0 0.105727f
c_58473 XI0.XI0.XI7.ZN_NEG 0 0.106313f
c_58482 XI0.XI0.XI10.ZN_NEG 0 0.105708f
c_58491 XI0.XI0.XI6.ZN_NEG 0 0.105776f
c_58501 XI0.XI0.XI9.ZN_NEG 0 0.105064f
c_58511 XI0.XI0.XI5.ZN_NEG 0 0.105802f
c_58519 XI0.XI0.XI8.ZN_NEG 0 0.108226f
c_58526 XI0.XI0.XI4.ZN_NEG 0 0.106004f
c_58541 XI0.XI1.XI4.XI3<0>.X 0 0.0735525f
c_58554 XI0.XI1.XI9.XI3<1>.Y 0 0.101377f
c_58568 XI0.XI1.XI15.XI3<0>.X 0 0.0750776f
c_58583 XI0.XI1.XI15.XI3<1>.Y 0 0.100391f
c_58596 XI0.XI1.XI4.XI3<1>.Y 0 0.100947f
c_58611 XI0.XI1.XI5.XI3<0>.X 0 0.0753132f
c_58624 XI0.XI1.XI5.XI3<1>.Y 0 0.100947f
c_58639 XI0.XI1.XI9.XI3<0>.X 0 0.0753187f
c_58654 XI0.XI1.XI8.XI3<0>.X 0 0.0752909f
c_58668 XI0.XI1.XI8.XI3<1>.Y 0 0.100943f
c_58682 XI0.XI1.XI12.XI3<0>.X 0 0.0753183f
c_58696 XI0.XI1.XI12.XI3<1>.Y 0 0.100947f
c_58710 XI0.XI1.XI13.XI3<0>.X 0 0.075316f
c_58724 XI0.XI1.XI13.XI3<1>.Y 0 0.100947f
c_58738 XI0.XI1.XI15.XI3<4>.X 0 0.0751318f
c_58753 XI0.XI1.XI15.XI3<5>.Y 0 0.101169f
c_58767 XI0.XI1.XI15.XI3<8>.X 0 0.0751344f
c_58784 XI0.XI1.XI15.XI3<9>.Y 0 0.100954f
c_58801 XI0.XI1.XI15.XI3<12>.X 0 0.0724775f
c_58819 XI0.XI1.XI15.XI3<13>.Y 0 0.0995373f
c_58833 XI0.XI1.XI15.XI3<2>.X 0 0.0796142f
c_58847 XI0.XI1.XI15.XI3<3>.Y 0 0.103078f
c_58860 XI0.XI1.XI15.XI3<3>.X 0 0.0782874f
c_58874 XI0.XI1.XI15.XI3<2>.Y 0 0.101965f
c_58888 XI0.XI1.XI15.XI3<3>.NEN 0 0.106176f
c_58902 XI0.XI1.XI15.XI3<2>.NEN 0 0.107094f
c_58915 XI0.XI1.XI15.XI3<1>.X 0 0.0749559f
c_58929 XI0.XI1.XI15.XI3<0>.Y 0 0.101434f
c_58944 XI0.XI1.XI15.XI3<1>.NEN 0 0.106171f
c_58958 XI0.XI1.XI15.XI3<0>.NEN 0 0.107707f
c_58972 XI0.XI1.XI15.XI3<6>.X 0 0.0746638f
c_58988 XI0.XI1.XI15.XI3<7>.Y 0 0.101034f
c_59002 XI0.XI1.XI15.XI3<7>.X 0 0.0748899f
c_59018 XI0.XI1.XI15.XI3<6>.Y 0 0.100481f
c_59033 XI0.XI1.XI15.XI3<7>.NEN 0 0.106268f
c_59049 XI0.XI1.XI15.XI3<6>.NEN 0 0.106996f
c_59062 XI0.XI1.XI15.XI3<5>.X 0 0.0749035f
c_59077 XI0.XI1.XI15.XI3<4>.Y 0 0.100023f
c_59092 XI0.XI1.XI15.XI3<5>.NEN 0 0.106171f
c_59107 XI0.XI1.XI15.XI3<4>.NEN 0 0.107094f
c_59123 XI0.XI1.XI15.XI3<10>.X 0 0.0746524f
c_59140 XI0.XI1.XI15.XI3<11>.Y 0 0.100488f
c_59155 XI0.XI1.XI15.XI3<11>.X 0 0.0746964f
c_59172 XI0.XI1.XI15.XI3<10>.Y 0 0.100459f
c_59188 XI0.XI1.XI15.XI3<11>.NEN 0 0.106331f
c_59203 XI0.XI1.XI15.XI3<10>.NEN 0 0.107207f
c_59217 XI0.XI1.XI15.XI3<9>.X 0 0.0753634f
c_59233 XI0.XI1.XI15.XI3<8>.Y 0 0.100452f
c_59249 XI0.XI1.XI15.XI3<9>.NEN 0 0.106181f
c_59265 XI0.XI1.XI15.XI3<8>.NEN 0 0.107094f
c_59283 XI0.XI1.XI15.XI3<14>.X 0 0.0718429f
c_59302 XI0.XI1.XI15.XI3<15>.Y 0 0.0991131f
c_59319 XI0.XI1.XI15.XI3<15>.X 0 0.0730439f
c_59339 XI0.XI1.XI15.XI3<14>.Y 0 0.0999451f
c_59353 XI0.XI1.XI15.XI3<15>.NEN 0 0.106783f
c_59369 XI0.XI1.XI15.XI3<14>.NEN 0 0.107105f
c_59384 XI0.XI1.XI15.XI3<13>.X 0 0.0734524f
c_59403 XI0.XI1.XI15.XI3<12>.Y 0 0.100417f
c_59419 XI0.XI1.XI15.XI3<13>.NEN 0 0.106174f
c_59435 XI0.XI1.XI15.XI3<12>.NEN 0 0.107119f
c_59447 XI0.XI1.XI3.XI3<0>.X 0 0.0759322f
c_59460 XI0.XI1.XI3.XI3<1>.Y 0 0.102068f
c_59474 XI0.XI1.XI3.XI3<4>.X 0 0.0741967f
c_59488 XI0.XI1.XI3.XI3<5>.Y 0 0.102197f
c_59502 XI0.XI1.XI3.XI3<8>.X 0 0.0742958f
c_59518 XI0.XI1.XI3.XI3<9>.Y 0 0.102298f
c_59533 XI0.XI1.XI3.XI3<12>.X 0 0.072483f
c_59550 XI0.XI1.XI3.XI3<13>.Y 0 0.100574f
c_59563 XI0.XI1.XI3.XI3<2>.X 0 0.0749299f
c_59576 XI0.XI1.XI3.XI3<3>.Y 0 0.101479f
c_59589 XI0.XI1.XI3.XI3<3>.X 0 0.0744642f
c_59603 XI0.XI1.XI3.XI3<2>.Y 0 0.10024f
c_59621 XI0.XI1.XI3.XI3<3>.NEN 0 0.0868961f
c_59639 XI0.XI1.XI3.XI3<2>.NEN 0 0.0875193f
c_59651 XI0.XI1.XI3.XI3<1>.X 0 0.075491f
c_59662 XI0.XI1.XI3.XI3<0>.Y 0 0.102656f
c_59680 XI0.XI1.XI3.XI3<1>.NEN 0 0.0868257f
c_59696 XI0.XI1.XI3.XI3<0>.NEN 0 0.0880916f
c_59710 XI0.XI1.XI3.XI3<6>.X 0 0.0725695f
c_59725 XI0.XI1.XI3.XI3<7>.Y 0 0.102035f
c_59739 XI0.XI1.XI3.XI3<7>.X 0 0.0730278f
c_59754 XI0.XI1.XI3.XI3<6>.Y 0 0.101386f
c_59773 XI0.XI1.XI3.XI3<7>.NEN 0 0.0869923f
c_59791 XI0.XI1.XI3.XI3<6>.NEN 0 0.0876548f
c_59804 XI0.XI1.XI3.XI3<5>.X 0 0.0746321f
c_59818 XI0.XI1.XI3.XI3<4>.Y 0 0.100409f
c_59837 XI0.XI1.XI3.XI3<5>.NEN 0 0.086949f
c_59856 XI0.XI1.XI3.XI3<4>.NEN 0 0.0876263f
c_59871 XI0.XI1.XI3.XI3<10>.X 0 0.0750129f
c_59887 XI0.XI1.XI3.XI3<11>.Y 0 0.101556f
c_59901 XI0.XI1.XI3.XI3<11>.X 0 0.0743077f
c_59917 XI0.XI1.XI3.XI3<10>.Y 0 0.100781f
c_59936 XI0.XI1.XI3.XI3<11>.NEN 0 0.0871811f
c_59955 XI0.XI1.XI3.XI3<10>.NEN 0 0.0875662f
c_59969 XI0.XI1.XI3.XI3<9>.X 0 0.0749807f
c_59984 XI0.XI1.XI3.XI3<8>.Y 0 0.101368f
c_60002 XI0.XI1.XI3.XI3<9>.NEN 0 0.0871345f
c_60021 XI0.XI1.XI3.XI3<8>.NEN 0 0.0875624f
c_60037 XI0.XI1.XI3.XI3<14>.X 0 0.0718695f
c_60054 XI0.XI1.XI3.XI3<15>.Y 0 0.0998181f
c_60070 XI0.XI1.XI3.XI3<15>.X 0 0.072612f
c_60088 XI0.XI1.XI3.XI3<14>.Y 0 0.100032f
c_60106 XI0.XI1.XI3.XI3<15>.NEN 0 0.0876455f
c_60126 XI0.XI1.XI3.XI3<14>.NEN 0 0.0876004f
c_60140 XI0.XI1.XI3.XI3<13>.X 0 0.0732749f
c_60157 XI0.XI1.XI3.XI3<12>.Y 0 0.100921f
c_60177 XI0.XI1.XI3.XI3<13>.NEN 0 0.0869494f
c_60196 XI0.XI1.XI3.XI3<12>.NEN 0 0.0877192f
c_60211 XI0.XI1.XI4.XI3<4>.X 0 0.0749138f
c_60226 XI0.XI1.XI4.XI3<5>.Y 0 0.101787f
c_60241 XI0.XI1.XI4.XI3<8>.X 0 0.0741974f
c_60258 XI0.XI1.XI4.XI3<9>.Y 0 0.101197f
c_60275 XI0.XI1.XI4.XI3<12>.X 0 0.0725462f
c_60293 XI0.XI1.XI4.XI3<13>.Y 0 0.100511f
c_60307 XI0.XI1.XI4.XI3<2>.X 0 0.0747644f
c_60321 XI0.XI1.XI4.XI3<3>.Y 0 0.100903f
c_60334 XI0.XI1.XI4.XI3<3>.X 0 0.074512f
c_60348 XI0.XI1.XI4.XI3<2>.Y 0 0.100281f
c_60366 XI0.XI1.XI4.XI3<3>.NEN 0 0.0868931f
c_60384 XI0.XI1.XI4.XI3<2>.NEN 0 0.0876294f
c_60397 XI0.XI1.XI4.XI3<1>.X 0 0.0750365f
c_60410 XI0.XI1.XI4.XI3<0>.Y 0 0.102155f
c_60427 XI0.XI1.XI4.XI3<1>.NEN 0 0.0868938f
c_60443 XI0.XI1.XI4.XI3<0>.NEN 0 0.0881863f
c_60457 XI0.XI1.XI4.XI3<6>.X 0 0.0750161f
c_60473 XI0.XI1.XI4.XI3<7>.Y 0 0.100957f
c_60488 XI0.XI1.XI4.XI3<7>.X 0 0.0745502f
c_60504 XI0.XI1.XI4.XI3<6>.Y 0 0.101068f
c_60522 XI0.XI1.XI4.XI3<7>.NEN 0 0.0870956f
c_60541 XI0.XI1.XI4.XI3<6>.NEN 0 0.0875468f
c_60555 XI0.XI1.XI4.XI3<5>.X 0 0.0728477f
c_60570 XI0.XI1.XI4.XI3<4>.Y 0 0.100211f
c_60588 XI0.XI1.XI4.XI3<5>.NEN 0 0.0870708f
c_60607 XI0.XI1.XI4.XI3<4>.NEN 0 0.0875051f
c_60623 XI0.XI1.XI4.XI3<10>.X 0 0.0745514f
c_60640 XI0.XI1.XI4.XI3<11>.Y 0 0.101408f
c_60655 XI0.XI1.XI4.XI3<11>.X 0 0.0748205f
c_60672 XI0.XI1.XI4.XI3<10>.Y 0 0.100591f
c_60690 XI0.XI1.XI4.XI3<11>.NEN 0 0.0872244f
c_60709 XI0.XI1.XI4.XI3<10>.NEN 0 0.0875864f
c_60724 XI0.XI1.XI4.XI3<9>.X 0 0.0745491f
c_60740 XI0.XI1.XI4.XI3<8>.Y 0 0.101177f
c_60759 XI0.XI1.XI4.XI3<9>.NEN 0 0.0869342f
c_60778 XI0.XI1.XI4.XI3<8>.NEN 0 0.0875468f
c_60795 XI0.XI1.XI4.XI3<14>.X 0 0.0725454f
c_60813 XI0.XI1.XI4.XI3<15>.Y 0 0.100086f
c_60830 XI0.XI1.XI4.XI3<15>.X 0 0.0735599f
c_60849 XI0.XI1.XI4.XI3<14>.Y 0 0.100725f
c_60867 XI0.XI1.XI4.XI3<15>.NEN 0 0.0876464f
c_60887 XI0.XI1.XI4.XI3<14>.NEN 0 0.0875701f
c_60903 XI0.XI1.XI4.XI3<13>.X 0 0.0736412f
c_60921 XI0.XI1.XI4.XI3<12>.Y 0 0.101311f
c_60941 XI0.XI1.XI4.XI3<13>.NEN 0 0.086943f
c_60960 XI0.XI1.XI4.XI3<12>.NEN 0 0.0877414f
c_60975 XI0.XI1.XI6.XI3<0>.X 0 0.075315f
c_60988 XI0.XI1.XI6.XI3<1>.Y 0 0.100947f
c_61002 XI0.XI1.XI6.XI3<4>.X 0 0.0747698f
c_61017 XI0.XI1.XI6.XI3<5>.Y 0 0.10152f
c_61032 XI0.XI1.XI6.XI3<8>.X 0 0.0748546f
c_61048 XI0.XI1.XI6.XI3<9>.Y 0 0.101356f
c_61065 XI0.XI1.XI6.XI3<12>.X 0 0.07287f
c_61083 XI0.XI1.XI6.XI3<13>.Y 0 0.100511f
c_61097 XI0.XI1.XI6.XI3<2>.X 0 0.0750422f
c_61111 XI0.XI1.XI6.XI3<3>.Y 0 0.100901f
c_61124 XI0.XI1.XI6.XI3<3>.X 0 0.0745673f
c_61138 XI0.XI1.XI6.XI3<2>.Y 0 0.100306f
c_61156 XI0.XI1.XI6.XI3<3>.NEN 0 0.0868931f
c_61174 XI0.XI1.XI6.XI3<2>.NEN 0 0.0876294f
c_61187 XI0.XI1.XI6.XI3<1>.X 0 0.0750372f
c_61200 XI0.XI1.XI6.XI3<0>.Y 0 0.102164f
c_61217 XI0.XI1.XI6.XI3<1>.NEN 0 0.0868938f
c_61233 XI0.XI1.XI6.XI3<0>.NEN 0 0.0882254f
c_61247 XI0.XI1.XI6.XI3<6>.X 0 0.0752697f
c_61263 XI0.XI1.XI6.XI3<7>.Y 0 0.101434f
c_61278 XI0.XI1.XI6.XI3<7>.X 0 0.0749457f
c_61293 XI0.XI1.XI6.XI3<6>.Y 0 0.101231f
c_61311 XI0.XI1.XI6.XI3<7>.NEN 0 0.0871095f
c_61330 XI0.XI1.XI6.XI3<6>.NEN 0 0.0875468f
c_61344 XI0.XI1.XI6.XI3<5>.X 0 0.0749434f
c_61359 XI0.XI1.XI6.XI3<4>.Y 0 0.100212f
c_61377 XI0.XI1.XI6.XI3<5>.NEN 0 0.087056f
c_61396 XI0.XI1.XI6.XI3<4>.NEN 0 0.0874208f
c_61412 XI0.XI1.XI6.XI3<10>.X 0 0.0748381f
c_61429 XI0.XI1.XI6.XI3<11>.Y 0 0.100952f
c_61444 XI0.XI1.XI6.XI3<11>.X 0 0.0748016f
c_61461 XI0.XI1.XI6.XI3<10>.Y 0 0.10059f
c_61480 XI0.XI1.XI6.XI3<11>.NEN 0 0.0871728f
c_61499 XI0.XI1.XI6.XI3<10>.NEN 0 0.0875864f
c_61514 XI0.XI1.XI6.XI3<9>.X 0 0.0745574f
c_61530 XI0.XI1.XI6.XI3<8>.Y 0 0.101236f
c_61549 XI0.XI1.XI6.XI3<9>.NEN 0 0.0869342f
c_61568 XI0.XI1.XI6.XI3<8>.NEN 0 0.087563f
c_61585 XI0.XI1.XI6.XI3<14>.X 0 0.0723887f
c_61603 XI0.XI1.XI6.XI3<15>.Y 0 0.100086f
c_61620 XI0.XI1.XI6.XI3<15>.X 0 0.0735654f
c_61639 XI0.XI1.XI6.XI3<14>.Y 0 0.100565f
c_61657 XI0.XI1.XI6.XI3<15>.NEN 0 0.0876766f
c_61677 XI0.XI1.XI6.XI3<14>.NEN 0 0.0875701f
c_61693 XI0.XI1.XI6.XI3<13>.X 0 0.0736484f
c_61711 XI0.XI1.XI6.XI3<12>.Y 0 0.101311f
c_61731 XI0.XI1.XI6.XI3<13>.NEN 0 0.086943f
c_61750 XI0.XI1.XI6.XI3<12>.NEN 0 0.0877414f
c_61764 XI0.XI1.XI5.XI3<4>.X 0 0.0747648f
c_61779 XI0.XI1.XI5.XI3<5>.Y 0 0.10152f
c_61794 XI0.XI1.XI5.XI3<8>.X 0 0.0748546f
c_61810 XI0.XI1.XI5.XI3<9>.Y 0 0.101356f
c_61826 XI0.XI1.XI5.XI3<12>.X 0 0.0728928f
c_61844 XI0.XI1.XI5.XI3<13>.Y 0 0.100511f
c_61858 XI0.XI1.XI5.XI3<2>.X 0 0.0785812f
c_61872 XI0.XI1.XI5.XI3<3>.Y 0 0.101098f
c_61885 XI0.XI1.XI5.XI3<3>.X 0 0.0756793f
c_61899 XI0.XI1.XI5.XI3<2>.Y 0 0.102053f
c_61917 XI0.XI1.XI5.XI3<3>.NEN 0 0.0868931f
c_61935 XI0.XI1.XI5.XI3<2>.NEN 0 0.0876223f
c_61948 XI0.XI1.XI5.XI3<1>.X 0 0.0749568f
c_61962 XI0.XI1.XI5.XI3<0>.Y 0 0.101991f
c_61979 XI0.XI1.XI5.XI3<1>.NEN 0 0.0868938f
c_61996 XI0.XI1.XI5.XI3<0>.NEN 0 0.0881404f
c_62010 XI0.XI1.XI5.XI3<6>.X 0 0.0752697f
c_62026 XI0.XI1.XI5.XI3<7>.Y 0 0.101401f
c_62041 XI0.XI1.XI5.XI3<7>.X 0 0.0749457f
c_62056 XI0.XI1.XI5.XI3<6>.Y 0 0.101231f
c_62074 XI0.XI1.XI5.XI3<7>.NEN 0 0.0871095f
c_62093 XI0.XI1.XI5.XI3<6>.NEN 0 0.0875468f
c_62107 XI0.XI1.XI5.XI3<5>.X 0 0.0749434f
c_62122 XI0.XI1.XI5.XI3<4>.Y 0 0.100214f
c_62140 XI0.XI1.XI5.XI3<5>.NEN 0 0.087056f
c_62158 XI0.XI1.XI5.XI3<4>.NEN 0 0.0875193f
c_62174 XI0.XI1.XI5.XI3<10>.X 0 0.0748381f
c_62191 XI0.XI1.XI5.XI3<11>.Y 0 0.101303f
c_62206 XI0.XI1.XI5.XI3<11>.X 0 0.0748016f
c_62223 XI0.XI1.XI5.XI3<10>.Y 0 0.100589f
c_62242 XI0.XI1.XI5.XI3<11>.NEN 0 0.0871719f
c_62261 XI0.XI1.XI5.XI3<10>.NEN 0 0.0875864f
c_62276 XI0.XI1.XI5.XI3<9>.X 0 0.0745574f
c_62292 XI0.XI1.XI5.XI3<8>.Y 0 0.101236f
c_62311 XI0.XI1.XI5.XI3<9>.NEN 0 0.0869342f
c_62330 XI0.XI1.XI5.XI3<8>.NEN 0 0.0875767f
c_62347 XI0.XI1.XI5.XI3<14>.X 0 0.0723887f
c_62365 XI0.XI1.XI5.XI3<15>.Y 0 0.100004f
c_62382 XI0.XI1.XI5.XI3<15>.X 0 0.073566f
c_62400 XI0.XI1.XI5.XI3<14>.Y 0 0.100728f
c_62418 XI0.XI1.XI5.XI3<15>.NEN 0 0.0876716f
c_62438 XI0.XI1.XI5.XI3<14>.NEN 0 0.0875701f
c_62454 XI0.XI1.XI5.XI3<13>.X 0 0.0736484f
c_62472 XI0.XI1.XI5.XI3<12>.Y 0 0.101311f
c_62492 XI0.XI1.XI5.XI3<13>.NEN 0 0.086947f
c_62511 XI0.XI1.XI5.XI3<12>.NEN 0 0.0877414f
c_62526 XI0.XI1.XI10.XI3<0>.X 0 0.0753166f
c_62539 XI0.XI1.XI10.XI3<1>.Y 0 0.100839f
c_62553 XI0.XI1.XI10.XI3<4>.X 0 0.0747648f
c_62568 XI0.XI1.XI10.XI3<5>.Y 0 0.101511f
c_62583 XI0.XI1.XI10.XI3<8>.X 0 0.0748546f
c_62599 XI0.XI1.XI10.XI3<9>.Y 0 0.10305f
c_62615 XI0.XI1.XI10.XI3<12>.X 0 0.0728928f
c_62633 XI0.XI1.XI10.XI3<13>.Y 0 0.100511f
c_62647 XI0.XI1.XI10.XI3<2>.X 0 0.0785692f
c_62661 XI0.XI1.XI10.XI3<3>.Y 0 0.100814f
c_62674 XI0.XI1.XI10.XI3<3>.X 0 0.0757948f
c_62688 XI0.XI1.XI10.XI3<2>.Y 0 0.102053f
c_62706 XI0.XI1.XI10.XI3<3>.NEN 0 0.0868951f
c_62724 XI0.XI1.XI10.XI3<2>.NEN 0 0.0875051f
c_62736 XI0.XI1.XI10.XI3<1>.X 0 0.0754703f
c_62750 XI0.XI1.XI10.XI3<0>.Y 0 0.102032f
c_62767 XI0.XI1.XI10.XI3<1>.NEN 0 0.0868938f
c_62784 XI0.XI1.XI10.XI3<0>.NEN 0 0.0882325f
c_62798 XI0.XI1.XI10.XI3<6>.X 0 0.0753324f
c_62814 XI0.XI1.XI10.XI3<7>.Y 0 0.101317f
c_62829 XI0.XI1.XI10.XI3<7>.X 0 0.0749457f
c_62844 XI0.XI1.XI10.XI3<6>.Y 0 0.10126f
c_62862 XI0.XI1.XI10.XI3<7>.NEN 0 0.0871095f
c_62881 XI0.XI1.XI10.XI3<6>.NEN 0 0.0875468f
c_62895 XI0.XI1.XI10.XI3<5>.X 0 0.07494f
c_62910 XI0.XI1.XI10.XI3<4>.Y 0 0.100058f
c_62928 XI0.XI1.XI10.XI3<5>.NEN 0 0.087056f
c_62946 XI0.XI1.XI10.XI3<4>.NEN 0 0.0875193f
c_62962 XI0.XI1.XI10.XI3<10>.X 0 0.0748381f
c_62979 XI0.XI1.XI10.XI3<11>.Y 0 0.101464f
c_62994 XI0.XI1.XI10.XI3<11>.X 0 0.0748016f
c_63011 XI0.XI1.XI10.XI3<10>.Y 0 0.100589f
c_63030 XI0.XI1.XI10.XI3<11>.NEN 0 0.0871714f
c_63049 XI0.XI1.XI10.XI3<10>.NEN 0 0.0875792f
c_63064 XI0.XI1.XI10.XI3<9>.X 0 0.0736655f
c_63080 XI0.XI1.XI10.XI3<8>.Y 0 0.101236f
c_63099 XI0.XI1.XI10.XI3<9>.NEN 0 0.0869529f
c_63118 XI0.XI1.XI10.XI3<8>.NEN 0 0.0875767f
c_63135 XI0.XI1.XI10.XI3<14>.X 0 0.0723887f
c_63153 XI0.XI1.XI10.XI3<15>.Y 0 0.0999863f
c_63170 XI0.XI1.XI10.XI3<15>.X 0 0.0735666f
c_63188 XI0.XI1.XI10.XI3<14>.Y 0 0.100728f
c_63206 XI0.XI1.XI10.XI3<15>.NEN 0 0.0876091f
c_63226 XI0.XI1.XI10.XI3<14>.NEN 0 0.0875701f
c_63243 XI0.XI1.XI10.XI3<13>.X 0 0.073538f
c_63261 XI0.XI1.XI10.XI3<12>.Y 0 0.101308f
c_63281 XI0.XI1.XI10.XI3<13>.NEN 0 0.086947f
c_63300 XI0.XI1.XI10.XI3<12>.NEN 0 0.087729f
c_63314 XI0.XI1.XI9.XI3<4>.X 0 0.0752609f
c_63329 XI0.XI1.XI9.XI3<5>.Y 0 0.101477f
c_63344 XI0.XI1.XI9.XI3<8>.X 0 0.0748546f
c_63360 XI0.XI1.XI9.XI3<9>.Y 0 0.103525f
c_63376 XI0.XI1.XI9.XI3<12>.X 0 0.0728928f
c_63394 XI0.XI1.XI9.XI3<13>.Y 0 0.100502f
c_63407 XI0.XI1.XI9.XI3<2>.X 0 0.0784206f
c_63421 XI0.XI1.XI9.XI3<3>.Y 0 0.100812f
c_63434 XI0.XI1.XI9.XI3<3>.X 0 0.0758441f
c_63448 XI0.XI1.XI9.XI3<2>.Y 0 0.102053f
c_63466 XI0.XI1.XI9.XI3<3>.NEN 0 0.0868992f
c_63484 XI0.XI1.XI9.XI3<2>.NEN 0 0.0874208f
c_63496 XI0.XI1.XI9.XI3<1>.X 0 0.0751195f
c_63510 XI0.XI1.XI9.XI3<0>.Y 0 0.102112f
c_63527 XI0.XI1.XI9.XI3<1>.NEN 0 0.0868938f
c_63544 XI0.XI1.XI9.XI3<0>.NEN 0 0.0881863f
c_63559 XI0.XI1.XI9.XI3<6>.X 0 0.0748347f
c_63574 XI0.XI1.XI9.XI3<7>.Y 0 0.101476f
c_63589 XI0.XI1.XI9.XI3<7>.X 0 0.0749491f
c_63604 XI0.XI1.XI9.XI3<6>.Y 0 0.101266f
c_63622 XI0.XI1.XI9.XI3<7>.NEN 0 0.0869906f
c_63641 XI0.XI1.XI9.XI3<6>.NEN 0 0.0875468f
c_63655 XI0.XI1.XI9.XI3<5>.X 0 0.07494f
c_63669 XI0.XI1.XI9.XI3<4>.Y 0 0.100218f
c_63687 XI0.XI1.XI9.XI3<5>.NEN 0 0.087001f
c_63705 XI0.XI1.XI9.XI3<4>.NEN 0 0.0875193f
c_63721 XI0.XI1.XI9.XI3<10>.X 0 0.0748381f
c_63738 XI0.XI1.XI9.XI3<11>.Y 0 0.101462f
c_63753 XI0.XI1.XI9.XI3<11>.X 0 0.0748016f
c_63770 XI0.XI1.XI9.XI3<10>.Y 0 0.10059f
c_63789 XI0.XI1.XI9.XI3<11>.NEN 0 0.0871733f
c_63808 XI0.XI1.XI9.XI3<10>.NEN 0 0.0875721f
c_63822 XI0.XI1.XI9.XI3<9>.X 0 0.0737546f
c_63838 XI0.XI1.XI9.XI3<8>.Y 0 0.101235f
c_63857 XI0.XI1.XI9.XI3<9>.NEN 0 0.0869859f
c_63876 XI0.XI1.XI9.XI3<8>.NEN 0 0.0875767f
c_63893 XI0.XI1.XI9.XI3<14>.X 0 0.0723887f
c_63911 XI0.XI1.XI9.XI3<15>.Y 0 0.0999109f
c_63928 XI0.XI1.XI9.XI3<15>.X 0 0.0735664f
c_63946 XI0.XI1.XI9.XI3<14>.Y 0 0.100728f
c_63964 XI0.XI1.XI9.XI3<15>.NEN 0 0.0875356f
c_63984 XI0.XI1.XI9.XI3<14>.NEN 0 0.0875701f
c_64000 XI0.XI1.XI9.XI3<13>.X 0 0.0738007f
c_64018 XI0.XI1.XI9.XI3<12>.Y 0 0.101148f
c_64038 XI0.XI1.XI9.XI3<13>.NEN 0 0.086947f
c_64057 XI0.XI1.XI9.XI3<12>.NEN 0 0.087729f
c_64072 XI0.XI1.XI7.XI3<0>.X 0 0.0753064f
c_64086 XI0.XI1.XI7.XI3<1>.Y 0 0.100762f
c_64100 XI0.XI1.XI7.XI3<4>.X 0 0.0752787f
c_64115 XI0.XI1.XI7.XI3<5>.Y 0 0.101353f
c_64130 XI0.XI1.XI7.XI3<8>.X 0 0.0748543f
c_64146 XI0.XI1.XI7.XI3<9>.Y 0 0.101959f
c_64162 XI0.XI1.XI7.XI3<12>.X 0 0.0728928f
c_64180 XI0.XI1.XI7.XI3<13>.Y 0 0.100469f
c_64193 XI0.XI1.XI7.XI3<2>.X 0 0.0784206f
c_64207 XI0.XI1.XI7.XI3<3>.Y 0 0.100813f
c_64221 XI0.XI1.XI7.XI3<3>.X 0 0.075737f
c_64235 XI0.XI1.XI7.XI3<2>.Y 0 0.102049f
c_64253 XI0.XI1.XI7.XI3<3>.NEN 0 0.0868992f
c_64270 XI0.XI1.XI7.XI3<2>.NEN 0 0.0875193f
c_64282 XI0.XI1.XI7.XI3<1>.X 0 0.0750456f
c_64296 XI0.XI1.XI7.XI3<0>.Y 0 0.102147f
c_64313 XI0.XI1.XI7.XI3<1>.NEN 0 0.0868938f
c_64330 XI0.XI1.XI7.XI3<0>.NEN 0 0.0881863f
c_64345 XI0.XI1.XI7.XI3<6>.X 0 0.0748347f
c_64360 XI0.XI1.XI7.XI3<7>.Y 0 0.101475f
c_64375 XI0.XI1.XI7.XI3<7>.X 0 0.0749491f
c_64390 XI0.XI1.XI7.XI3<6>.Y 0 0.101266f
c_64408 XI0.XI1.XI7.XI3<7>.NEN 0 0.0869906f
c_64427 XI0.XI1.XI7.XI3<6>.NEN 0 0.0875468f
c_64441 XI0.XI1.XI7.XI3<5>.X 0 0.0749998f
c_64455 XI0.XI1.XI7.XI3<4>.Y 0 0.100218f
c_64473 XI0.XI1.XI7.XI3<5>.NEN 0 0.0870009f
c_64491 XI0.XI1.XI7.XI3<4>.NEN 0 0.0875193f
c_64507 XI0.XI1.XI7.XI3<10>.X 0 0.0748233f
c_64524 XI0.XI1.XI7.XI3<11>.Y 0 0.101461f
c_64539 XI0.XI1.XI7.XI3<11>.X 0 0.0748016f
c_64556 XI0.XI1.XI7.XI3<10>.Y 0 0.10059f
c_64575 XI0.XI1.XI7.XI3<11>.NEN 0 0.0871905f
c_64594 XI0.XI1.XI7.XI3<10>.NEN 0 0.0874878f
c_64608 XI0.XI1.XI7.XI3<9>.X 0 0.0743231f
c_64624 XI0.XI1.XI7.XI3<8>.Y 0 0.101235f
c_64643 XI0.XI1.XI7.XI3<9>.NEN 0 0.0869859f
c_64662 XI0.XI1.XI7.XI3<8>.NEN 0 0.0875767f
c_64680 XI0.XI1.XI7.XI3<14>.X 0 0.0723887f
c_64697 XI0.XI1.XI7.XI3<15>.Y 0 0.100091f
c_64714 XI0.XI1.XI7.XI3<15>.X 0 0.0735657f
c_64732 XI0.XI1.XI7.XI3<14>.Y 0 0.100728f
c_64749 XI0.XI1.XI7.XI3<15>.NEN 0 0.0876798f
c_64769 XI0.XI1.XI7.XI3<14>.NEN 0 0.0875701f
c_64785 XI0.XI1.XI7.XI3<13>.X 0 0.0738007f
c_64802 XI0.XI1.XI7.XI3<12>.Y 0 0.101311f
c_64822 XI0.XI1.XI7.XI3<13>.NEN 0 0.086947f
c_64841 XI0.XI1.XI7.XI3<12>.NEN 0 0.087729f
c_64855 XI0.XI1.XI8.XI3<4>.X 0 0.0752991f
c_64870 XI0.XI1.XI8.XI3<5>.Y 0 0.101269f
c_64885 XI0.XI1.XI8.XI3<8>.X 0 0.0748437f
c_64901 XI0.XI1.XI8.XI3<9>.Y 0 0.101963f
c_64917 XI0.XI1.XI8.XI3<12>.X 0 0.0728928f
c_64935 XI0.XI1.XI8.XI3<13>.Y 0 0.100437f
c_64948 XI0.XI1.XI8.XI3<2>.X 0 0.0784206f
c_64962 XI0.XI1.XI8.XI3<3>.Y 0 0.100804f
c_64975 XI0.XI1.XI8.XI3<3>.X 0 0.0769124f
c_64989 XI0.XI1.XI8.XI3<2>.Y 0 0.101895f
c_65007 XI0.XI1.XI8.XI3<3>.NEN 0 0.0868992f
c_65024 XI0.XI1.XI8.XI3<2>.NEN 0 0.0875193f
c_65036 XI0.XI1.XI8.XI3<1>.X 0 0.0750456f
c_65050 XI0.XI1.XI8.XI3<0>.Y 0 0.102198f
c_65067 XI0.XI1.XI8.XI3<1>.NEN 0 0.0868938f
c_65084 XI0.XI1.XI8.XI3<0>.NEN 0 0.0882353f
c_65099 XI0.XI1.XI8.XI3<6>.X 0 0.0748347f
c_65114 XI0.XI1.XI8.XI3<7>.Y 0 0.101475f
c_65129 XI0.XI1.XI8.XI3<7>.X 0 0.07486f
c_65144 XI0.XI1.XI8.XI3<6>.Y 0 0.101266f
c_65162 XI0.XI1.XI8.XI3<7>.NEN 0 0.0869906f
c_65181 XI0.XI1.XI8.XI3<6>.NEN 0 0.0875468f
c_65195 XI0.XI1.XI8.XI3<5>.X 0 0.0749998f
c_65209 XI0.XI1.XI8.XI3<4>.Y 0 0.100243f
c_65227 XI0.XI1.XI8.XI3<5>.NEN 0 0.0870009f
c_65245 XI0.XI1.XI8.XI3<4>.NEN 0 0.0875193f
c_65261 XI0.XI1.XI8.XI3<10>.X 0 0.0748233f
c_65278 XI0.XI1.XI8.XI3<11>.Y 0 0.101462f
c_65293 XI0.XI1.XI8.XI3<11>.X 0 0.0748016f
c_65310 XI0.XI1.XI8.XI3<10>.Y 0 0.100586f
c_65329 XI0.XI1.XI8.XI3<11>.NEN 0 0.0871762f
c_65347 XI0.XI1.XI8.XI3<10>.NEN 0 0.0875864f
c_65361 XI0.XI1.XI8.XI3<9>.X 0 0.0750082f
c_65377 XI0.XI1.XI8.XI3<8>.Y 0 0.101235f
c_65396 XI0.XI1.XI8.XI3<9>.NEN 0 0.0869859f
c_65415 XI0.XI1.XI8.XI3<8>.NEN 0 0.0875767f
c_65433 XI0.XI1.XI8.XI3<14>.X 0 0.0723887f
c_65450 XI0.XI1.XI8.XI3<15>.Y 0 0.100119f
c_65467 XI0.XI1.XI8.XI3<15>.X 0 0.0735656f
c_65485 XI0.XI1.XI8.XI3<14>.Y 0 0.100728f
c_65502 XI0.XI1.XI8.XI3<15>.NEN 0 0.0876589f
c_65522 XI0.XI1.XI8.XI3<14>.NEN 0 0.0875701f
c_65538 XI0.XI1.XI8.XI3<13>.X 0 0.0738007f
c_65555 XI0.XI1.XI8.XI3<12>.Y 0 0.101311f
c_65575 XI0.XI1.XI8.XI3<13>.NEN 0 0.086947f
c_65594 XI0.XI1.XI8.XI3<12>.NEN 0 0.087729f
c_65608 XI0.XI1.XI11.XI3<0>.X 0 0.0753144f
c_65622 XI0.XI1.XI11.XI3<1>.Y 0 0.100947f
c_65636 XI0.XI1.XI11.XI3<4>.X 0 0.0752871f
c_65650 XI0.XI1.XI11.XI3<5>.Y 0 0.10152f
c_65665 XI0.XI1.XI11.XI3<8>.X 0 0.0748317f
c_65681 XI0.XI1.XI11.XI3<9>.Y 0 0.101963f
c_65697 XI0.XI1.XI11.XI3<12>.X 0 0.0728928f
c_65715 XI0.XI1.XI11.XI3<13>.Y 0 0.10035f
c_65728 XI0.XI1.XI11.XI3<2>.X 0 0.0784206f
c_65742 XI0.XI1.XI11.XI3<3>.Y 0 0.102987f
c_65755 XI0.XI1.XI11.XI3<3>.X 0 0.076201f
c_65768 XI0.XI1.XI11.XI3<2>.Y 0 0.102053f
c_65786 XI0.XI1.XI11.XI3<3>.NEN 0 0.0868992f
c_65803 XI0.XI1.XI11.XI3<2>.NEN 0 0.0875193f
c_65815 XI0.XI1.XI11.XI3<1>.X 0 0.0750456f
c_65829 XI0.XI1.XI11.XI3<0>.Y 0 0.10221f
c_65847 XI0.XI1.XI11.XI3<1>.NEN 0 0.0867791f
c_65865 XI0.XI1.XI11.XI3<0>.NEN 0 0.0879949f
c_65880 XI0.XI1.XI11.XI3<6>.X 0 0.0748347f
c_65895 XI0.XI1.XI11.XI3<7>.Y 0 0.101475f
c_65909 XI0.XI1.XI11.XI3<7>.X 0 0.0749491f
c_65924 XI0.XI1.XI11.XI3<6>.Y 0 0.101266f
c_65942 XI0.XI1.XI11.XI3<7>.NEN 0 0.0870011f
c_65961 XI0.XI1.XI11.XI3<6>.NEN 0 0.0875468f
c_65975 XI0.XI1.XI11.XI3<5>.X 0 0.0749362f
c_65989 XI0.XI1.XI11.XI3<4>.Y 0 0.10028f
c_66007 XI0.XI1.XI11.XI3<5>.NEN 0 0.0868938f
c_66025 XI0.XI1.XI11.XI3<4>.NEN 0 0.0875193f
c_66041 XI0.XI1.XI11.XI3<10>.X 0 0.0748233f
c_66058 XI0.XI1.XI11.XI3<11>.Y 0 0.101909f
c_66073 XI0.XI1.XI11.XI3<11>.X 0 0.0748016f
c_66090 XI0.XI1.XI11.XI3<10>.Y 0 0.100425f
c_66109 XI0.XI1.XI11.XI3<11>.NEN 0 0.0871757f
c_66127 XI0.XI1.XI11.XI3<10>.NEN 0 0.0875864f
c_66141 XI0.XI1.XI11.XI3<9>.X 0 0.0750237f
c_66157 XI0.XI1.XI11.XI3<8>.Y 0 0.101235f
c_66176 XI0.XI1.XI11.XI3<9>.NEN 0 0.0869859f
c_66195 XI0.XI1.XI11.XI3<8>.NEN 0 0.0875767f
c_66213 XI0.XI1.XI11.XI3<14>.X 0 0.0723887f
c_66230 XI0.XI1.XI11.XI3<15>.Y 0 0.100048f
c_66247 XI0.XI1.XI11.XI3<15>.X 0 0.0735663f
c_66266 XI0.XI1.XI11.XI3<14>.Y 0 0.100541f
c_66283 XI0.XI1.XI11.XI3<15>.NEN 0 0.0877016f
c_66303 XI0.XI1.XI11.XI3<14>.NEN 0 0.0875826f
c_66319 XI0.XI1.XI11.XI3<13>.X 0 0.0738007f
c_66336 XI0.XI1.XI11.XI3<12>.Y 0 0.101311f
c_66356 XI0.XI1.XI11.XI3<13>.NEN 0 0.0869449f
c_66375 XI0.XI1.XI11.XI3<12>.NEN 0 0.087729f
c_66389 XI0.XI1.XI12.XI3<4>.X 0 0.0752871f
c_66403 XI0.XI1.XI12.XI3<5>.Y 0 0.101519f
c_66417 XI0.XI1.XI12.XI3<8>.X 0 0.0748546f
c_66433 XI0.XI1.XI12.XI3<9>.Y 0 0.101963f
c_66450 XI0.XI1.XI12.XI3<12>.X 0 0.0728928f
c_66467 XI0.XI1.XI12.XI3<13>.Y 0 0.100511f
c_66480 XI0.XI1.XI12.XI3<2>.X 0 0.0784256f
c_66494 XI0.XI1.XI12.XI3<3>.Y 0 0.102955f
c_66507 XI0.XI1.XI12.XI3<3>.X 0 0.0765056f
c_66520 XI0.XI1.XI12.XI3<2>.Y 0 0.10246f
c_66538 XI0.XI1.XI12.XI3<3>.NEN 0 0.0868992f
c_66555 XI0.XI1.XI12.XI3<2>.NEN 0 0.0875193f
c_66568 XI0.XI1.XI12.XI3<1>.X 0 0.0749419f
c_66582 XI0.XI1.XI12.XI3<0>.Y 0 0.102175f
c_66600 XI0.XI1.XI12.XI3<1>.NEN 0 0.0868526f
c_66617 XI0.XI1.XI12.XI3<0>.NEN 0 0.0881263f
c_66632 XI0.XI1.XI12.XI3<6>.X 0 0.0748347f
c_66647 XI0.XI1.XI12.XI3<7>.Y 0 0.101552f
c_66661 XI0.XI1.XI12.XI3<7>.X 0 0.0749491f
c_66676 XI0.XI1.XI12.XI3<6>.Y 0 0.101265f
c_66694 XI0.XI1.XI12.XI3<7>.NEN 0 0.0870022f
c_66713 XI0.XI1.XI12.XI3<6>.NEN 0 0.0875468f
c_66727 XI0.XI1.XI12.XI3<5>.X 0 0.0749362f
c_66741 XI0.XI1.XI12.XI3<4>.Y 0 0.10028f
c_66759 XI0.XI1.XI12.XI3<5>.NEN 0 0.0868938f
c_66777 XI0.XI1.XI12.XI3<4>.NEN 0 0.0875193f
c_66793 XI0.XI1.XI12.XI3<10>.X 0 0.0748233f
c_66810 XI0.XI1.XI12.XI3<11>.Y 0 0.101876f
c_66825 XI0.XI1.XI12.XI3<11>.X 0 0.0748016f
c_66841 XI0.XI1.XI12.XI3<10>.Y 0 0.100588f
c_66860 XI0.XI1.XI12.XI3<11>.NEN 0 0.0871742f
c_66878 XI0.XI1.XI12.XI3<10>.NEN 0 0.0875864f
c_66892 XI0.XI1.XI12.XI3<9>.X 0 0.0754565f
c_66908 XI0.XI1.XI12.XI3<8>.Y 0 0.101235f
c_66927 XI0.XI1.XI12.XI3<9>.NEN 0 0.0869866f
c_66946 XI0.XI1.XI12.XI3<8>.NEN 0 0.0875767f
c_66964 XI0.XI1.XI12.XI3<14>.X 0 0.0723887f
c_66981 XI0.XI1.XI12.XI3<15>.Y 0 0.100064f
c_66998 XI0.XI1.XI12.XI3<15>.X 0 0.0735248f
c_67017 XI0.XI1.XI12.XI3<14>.Y 0 0.100617f
c_67034 XI0.XI1.XI12.XI3<15>.NEN 0 0.0876148f
c_67054 XI0.XI1.XI12.XI3<14>.NEN 0 0.0875826f
c_67070 XI0.XI1.XI12.XI3<13>.X 0 0.0738007f
c_67087 XI0.XI1.XI12.XI3<12>.Y 0 0.101311f
c_67107 XI0.XI1.XI12.XI3<13>.NEN 0 0.0869356f
c_67126 XI0.XI1.XI12.XI3<12>.NEN 0 0.087729f
c_67140 XI0.XI1.XI14.XI3<0>.X 0 0.0753192f
c_67154 XI0.XI1.XI14.XI3<1>.Y 0 0.100947f
c_67168 XI0.XI1.XI14.XI3<4>.X 0 0.0752871f
c_67182 XI0.XI1.XI14.XI3<5>.Y 0 0.10152f
c_67196 XI0.XI1.XI14.XI3<8>.X 0 0.0748546f
c_67212 XI0.XI1.XI14.XI3<9>.Y 0 0.101963f
c_67229 XI0.XI1.XI14.XI3<12>.X 0 0.0728928f
c_67246 XI0.XI1.XI14.XI3<13>.Y 0 0.100511f
c_67259 XI0.XI1.XI14.XI3<2>.X 0 0.0747644f
c_67273 XI0.XI1.XI14.XI3<3>.Y 0 0.102872f
c_67287 XI0.XI1.XI14.XI3<3>.X 0 0.07528f
c_67300 XI0.XI1.XI14.XI3<2>.Y 0 0.100281f
c_67318 XI0.XI1.XI14.XI3<3>.NEN 0 0.0868257f
c_67335 XI0.XI1.XI14.XI3<2>.NEN 0 0.0875193f
c_67348 XI0.XI1.XI14.XI3<1>.X 0 0.0750284f
c_67362 XI0.XI1.XI14.XI3<0>.Y 0 0.102034f
c_67380 XI0.XI1.XI14.XI3<1>.NEN 0 0.086883f
c_67397 XI0.XI1.XI14.XI3<0>.NEN 0 0.0880698f
c_67412 XI0.XI1.XI14.XI3<6>.X 0 0.0748238f
c_67427 XI0.XI1.XI14.XI3<7>.Y 0 0.10158f
c_67441 XI0.XI1.XI14.XI3<7>.X 0 0.0749491f
c_67456 XI0.XI1.XI14.XI3<6>.Y 0 0.101266f
c_67474 XI0.XI1.XI14.XI3<7>.NEN 0 0.0870033f
c_67493 XI0.XI1.XI14.XI3<6>.NEN 0 0.0875397f
c_67507 XI0.XI1.XI14.XI3<5>.X 0 0.0748471f
c_67522 XI0.XI1.XI14.XI3<4>.Y 0 0.100097f
c_67540 XI0.XI1.XI14.XI3<5>.NEN 0 0.0868938f
c_67558 XI0.XI1.XI14.XI3<4>.NEN 0 0.0875193f
c_67574 XI0.XI1.XI14.XI3<10>.X 0 0.0748233f
c_67591 XI0.XI1.XI14.XI3<11>.Y 0 0.101387f
c_67606 XI0.XI1.XI14.XI3<11>.X 0 0.0748016f
c_67622 XI0.XI1.XI14.XI3<10>.Y 0 0.100588f
c_67641 XI0.XI1.XI14.XI3<11>.NEN 0 0.0871723f
c_67659 XI0.XI1.XI14.XI3<10>.NEN 0 0.0875864f
c_67673 XI0.XI1.XI14.XI3<9>.X 0 0.0754565f
c_67689 XI0.XI1.XI14.XI3<8>.Y 0 0.101231f
c_67708 XI0.XI1.XI14.XI3<9>.NEN 0 0.0869866f
c_67727 XI0.XI1.XI14.XI3<8>.NEN 0 0.0875468f
c_67745 XI0.XI1.XI14.XI3<14>.X 0 0.0723887f
c_67762 XI0.XI1.XI14.XI3<15>.Y 0 0.100088f
c_67779 XI0.XI1.XI14.XI3<15>.X 0 0.0735244f
c_67798 XI0.XI1.XI14.XI3<14>.Y 0 0.100677f
c_67815 XI0.XI1.XI14.XI3<15>.NEN 0 0.0876091f
c_67835 XI0.XI1.XI14.XI3<14>.NEN 0 0.0875826f
c_67851 XI0.XI1.XI14.XI3<13>.X 0 0.0738007f
c_67868 XI0.XI1.XI14.XI3<12>.Y 0 0.101311f
c_67888 XI0.XI1.XI14.XI3<13>.NEN 0 0.0869356f
c_67907 XI0.XI1.XI14.XI3<12>.NEN 0 0.087729f
c_67921 XI0.XI1.XI13.XI3<4>.X 0 0.0752871f
c_67935 XI0.XI1.XI13.XI3<5>.Y 0 0.10152f
c_67949 XI0.XI1.XI13.XI3<8>.X 0 0.0748546f
c_67965 XI0.XI1.XI13.XI3<9>.Y 0 0.101955f
c_67982 XI0.XI1.XI13.XI3<12>.X 0 0.0728928f
c_67999 XI0.XI1.XI13.XI3<13>.Y 0 0.100511f
c_68013 XI0.XI1.XI13.XI3<2>.X 0 0.0784206f
c_68026 XI0.XI1.XI13.XI3<3>.Y 0 0.103171f
c_68039 XI0.XI1.XI13.XI3<3>.X 0 0.0780287f
c_68052 XI0.XI1.XI13.XI3<2>.Y 0 0.102053f
c_68069 XI0.XI1.XI13.XI3<3>.NEN 0 0.0868992f
c_68086 XI0.XI1.XI13.XI3<2>.NEN 0 0.0875193f
c_68099 XI0.XI1.XI13.XI3<1>.X 0 0.0750456f
c_68112 XI0.XI1.XI13.XI3<0>.Y 0 0.102194f
c_68130 XI0.XI1.XI13.XI3<1>.NEN 0 0.0868938f
c_68147 XI0.XI1.XI13.XI3<0>.NEN 0 0.0880683f
c_68162 XI0.XI1.XI13.XI3<6>.X 0 0.0748117f
c_68177 XI0.XI1.XI13.XI3<7>.Y 0 0.101574f
c_68191 XI0.XI1.XI13.XI3<7>.X 0 0.0749491f
c_68206 XI0.XI1.XI13.XI3<6>.Y 0 0.101266f
c_68224 XI0.XI1.XI13.XI3<7>.NEN 0 0.0870284f
c_68243 XI0.XI1.XI13.XI3<6>.NEN 0 0.0875326f
c_68256 XI0.XI1.XI13.XI3<5>.X 0 0.0749362f
c_68270 XI0.XI1.XI13.XI3<4>.Y 0 0.100334f
c_68288 XI0.XI1.XI13.XI3<5>.NEN 0 0.0868938f
c_68306 XI0.XI1.XI13.XI3<4>.NEN 0 0.0875193f
c_68322 XI0.XI1.XI13.XI3<10>.X 0 0.0748233f
c_68339 XI0.XI1.XI13.XI3<11>.Y 0 0.101302f
c_68354 XI0.XI1.XI13.XI3<11>.X 0 0.0748016f
c_68370 XI0.XI1.XI13.XI3<10>.Y 0 0.101242f
c_68389 XI0.XI1.XI13.XI3<11>.NEN 0 0.0871723f
c_68407 XI0.XI1.XI13.XI3<10>.NEN 0 0.0875864f
c_68421 XI0.XI1.XI13.XI3<9>.X 0 0.0754531f
c_68437 XI0.XI1.XI13.XI3<8>.Y 0 0.101071f
c_68456 XI0.XI1.XI13.XI3<9>.NEN 0 0.0869866f
c_68475 XI0.XI1.XI13.XI3<8>.NEN 0 0.0875468f
c_68493 XI0.XI1.XI13.XI3<14>.X 0 0.0723887f
c_68511 XI0.XI1.XI13.XI3<15>.Y 0 0.0999005f
c_68528 XI0.XI1.XI13.XI3<15>.X 0 0.0735237f
c_68547 XI0.XI1.XI13.XI3<14>.Y 0 0.100702f
c_68564 XI0.XI1.XI13.XI3<15>.NEN 0 0.0877089f
c_68584 XI0.XI1.XI13.XI3<14>.NEN 0 0.0875754f
c_68600 XI0.XI1.XI13.XI3<13>.X 0 0.0737014f
c_68618 XI0.XI1.XI13.XI3<12>.Y 0 0.101125f
c_68638 XI0.XI1.XI13.XI3<13>.NEN 0 0.0869316f
c_68657 XI0.XI1.XI13.XI3<12>.NEN 0 0.0877414f
c_68926 XI2.NET1<0> 0 4.43296f
c_69195 XI2.NET1<1> 0 4.40853f
c_69465 XI2.NET1<2> 0 4.44509f
c_69736 XI2.NET1<3> 0 4.48973f
c_70009 XI2.NET1<4> 0 4.49113f
c_70282 XI2.NET1<5> 0 4.49876f
c_70557 XI2.NET1<6> 0 4.5368f
c_70831 XI2.NET1<7> 0 4.53628f
c_71108 XI2.NET1<8> 0 4.58911f
c_71385 XI2.NET1<9> 0 4.6007f
c_71660 XI2.NET1<10> 0 4.53273f
c_71934 XI2.NET1<11> 0 4.66079f
c_72191 XI2.NET1<12> 0 4.7231f
c_72199 XI2.XI0.NET_11XX 0 0.15093f
c_72229 XI2.XI0.NET_XX00 0 1.10724f
c_72251 XI2.XI0.NET_XX11 0 0.70712f
c_72268 XI2.XI0.NET_10XX 0 0.637731f
c_72284 XI2.XI0.ADDR_BAR<2> 0 0.636229f
c_72301 XI2.XI0.ADDR_BAR<0> 0 0.70305f
c_72325 XI2.XI0.NET_XX10 0 0.981912f
c_72343 XI2.XI0.NET_01XX 0 0.614487f
c_72358 XI2.XI0.ADDR_BAR<1> 0 0.466041f
c_72379 XI2.XI0.NET_XX01 0 0.972175f
c_72396 XI2.XI0.NET_00XX 0 0.630231f
c_72413 XI2.XI0.ADDR_BAR<3> 0 0.381154f
c_72420 XI2.XI0.XI11.ZN_NEG 0 0.105727f
c_72428 XI2.XI0.XI7.ZN_NEG 0 0.106341f
c_72437 XI2.XI0.XI10.ZN_NEG 0 0.105718f
c_72446 XI2.XI0.XI6.ZN_NEG 0 0.105791f
c_72456 XI2.XI0.XI9.ZN_NEG 0 0.105064f
c_72466 XI2.XI0.XI5.ZN_NEG 0 0.105802f
c_72474 XI2.XI0.XI8.ZN_NEG 0 0.108226f
c_72481 XI2.XI0.XI4.ZN_NEG 0 0.106004f
c_72496 XI2.XI1.XI4.XI3<0>.X 0 0.0735525f
c_72509 XI2.XI1.XI9.XI3<1>.Y 0 0.101377f
c_72523 XI2.XI1.XI15.XI3<0>.X 0 0.0750776f
c_72538 XI2.XI1.XI15.XI3<1>.Y 0 0.100391f
c_72551 XI2.XI1.XI4.XI3<1>.Y 0 0.100947f
c_72566 XI2.XI1.XI5.XI3<0>.X 0 0.0753132f
c_72579 XI2.XI1.XI5.XI3<1>.Y 0 0.100947f
c_72594 XI2.XI1.XI9.XI3<0>.X 0 0.0753187f
c_72609 XI2.XI1.XI8.XI3<0>.X 0 0.0752909f
c_72623 XI2.XI1.XI8.XI3<1>.Y 0 0.100943f
c_72637 XI2.XI1.XI12.XI3<0>.X 0 0.0753183f
c_72651 XI2.XI1.XI12.XI3<1>.Y 0 0.100947f
c_72665 XI2.XI1.XI13.XI3<0>.X 0 0.075316f
c_72679 XI2.XI1.XI13.XI3<1>.Y 0 0.100947f
c_72693 XI2.XI1.XI15.XI3<4>.X 0 0.0751318f
c_72708 XI2.XI1.XI15.XI3<5>.Y 0 0.101169f
c_72722 XI2.XI1.XI15.XI3<8>.X 0 0.0751344f
c_72739 XI2.XI1.XI15.XI3<9>.Y 0 0.100954f
c_72756 XI2.XI1.XI15.XI3<12>.X 0 0.0724775f
c_72774 XI2.XI1.XI15.XI3<13>.Y 0 0.0995373f
c_72788 XI2.XI1.XI15.XI3<2>.X 0 0.0796142f
c_72802 XI2.XI1.XI15.XI3<3>.Y 0 0.103078f
c_72815 XI2.XI1.XI15.XI3<3>.X 0 0.0782874f
c_72829 XI2.XI1.XI15.XI3<2>.Y 0 0.101965f
c_72843 XI2.XI1.XI15.XI3<3>.NEN 0 0.106176f
c_72857 XI2.XI1.XI15.XI3<2>.NEN 0 0.107094f
c_72870 XI2.XI1.XI15.XI3<1>.X 0 0.0749559f
c_72884 XI2.XI1.XI15.XI3<0>.Y 0 0.101434f
c_72899 XI2.XI1.XI15.XI3<1>.NEN 0 0.106171f
c_72913 XI2.XI1.XI15.XI3<0>.NEN 0 0.107707f
c_72927 XI2.XI1.XI15.XI3<6>.X 0 0.0746638f
c_72943 XI2.XI1.XI15.XI3<7>.Y 0 0.101034f
c_72957 XI2.XI1.XI15.XI3<7>.X 0 0.0748899f
c_72973 XI2.XI1.XI15.XI3<6>.Y 0 0.100481f
c_72988 XI2.XI1.XI15.XI3<7>.NEN 0 0.106268f
c_73004 XI2.XI1.XI15.XI3<6>.NEN 0 0.106996f
c_73017 XI2.XI1.XI15.XI3<5>.X 0 0.0749035f
c_73032 XI2.XI1.XI15.XI3<4>.Y 0 0.100023f
c_73047 XI2.XI1.XI15.XI3<5>.NEN 0 0.106171f
c_73062 XI2.XI1.XI15.XI3<4>.NEN 0 0.107094f
c_73078 XI2.XI1.XI15.XI3<10>.X 0 0.0746524f
c_73095 XI2.XI1.XI15.XI3<11>.Y 0 0.100488f
c_73110 XI2.XI1.XI15.XI3<11>.X 0 0.0746964f
c_73127 XI2.XI1.XI15.XI3<10>.Y 0 0.100459f
c_73143 XI2.XI1.XI15.XI3<11>.NEN 0 0.106331f
c_73158 XI2.XI1.XI15.XI3<10>.NEN 0 0.107207f
c_73172 XI2.XI1.XI15.XI3<9>.X 0 0.0753634f
c_73188 XI2.XI1.XI15.XI3<8>.Y 0 0.100452f
c_73204 XI2.XI1.XI15.XI3<9>.NEN 0 0.106181f
c_73220 XI2.XI1.XI15.XI3<8>.NEN 0 0.107094f
c_73238 XI2.XI1.XI15.XI3<14>.X 0 0.0718429f
c_73257 XI2.XI1.XI15.XI3<15>.Y 0 0.0991131f
c_73274 XI2.XI1.XI15.XI3<15>.X 0 0.0730439f
c_73294 XI2.XI1.XI15.XI3<14>.Y 0 0.0999451f
c_73308 XI2.XI1.XI15.XI3<15>.NEN 0 0.106783f
c_73324 XI2.XI1.XI15.XI3<14>.NEN 0 0.107105f
c_73339 XI2.XI1.XI15.XI3<13>.X 0 0.0734524f
c_73358 XI2.XI1.XI15.XI3<12>.Y 0 0.100417f
c_73374 XI2.XI1.XI15.XI3<13>.NEN 0 0.106174f
c_73390 XI2.XI1.XI15.XI3<12>.NEN 0 0.107119f
c_73402 XI2.XI1.XI3.XI3<0>.X 0 0.0759322f
c_73415 XI2.XI1.XI3.XI3<1>.Y 0 0.102068f
c_73429 XI2.XI1.XI3.XI3<4>.X 0 0.0741967f
c_73443 XI2.XI1.XI3.XI3<5>.Y 0 0.102197f
c_73457 XI2.XI1.XI3.XI3<8>.X 0 0.0742958f
c_73473 XI2.XI1.XI3.XI3<9>.Y 0 0.102298f
c_73488 XI2.XI1.XI3.XI3<12>.X 0 0.072483f
c_73505 XI2.XI1.XI3.XI3<13>.Y 0 0.100574f
c_73518 XI2.XI1.XI3.XI3<2>.X 0 0.0749299f
c_73531 XI2.XI1.XI3.XI3<3>.Y 0 0.101479f
c_73544 XI2.XI1.XI3.XI3<3>.X 0 0.0744642f
c_73558 XI2.XI1.XI3.XI3<2>.Y 0 0.10024f
c_73576 XI2.XI1.XI3.XI3<3>.NEN 0 0.0868961f
c_73594 XI2.XI1.XI3.XI3<2>.NEN 0 0.0875193f
c_73606 XI2.XI1.XI3.XI3<1>.X 0 0.075491f
c_73617 XI2.XI1.XI3.XI3<0>.Y 0 0.102656f
c_73635 XI2.XI1.XI3.XI3<1>.NEN 0 0.0868257f
c_73651 XI2.XI1.XI3.XI3<0>.NEN 0 0.0880916f
c_73665 XI2.XI1.XI3.XI3<6>.X 0 0.0725695f
c_73680 XI2.XI1.XI3.XI3<7>.Y 0 0.102035f
c_73694 XI2.XI1.XI3.XI3<7>.X 0 0.0730278f
c_73709 XI2.XI1.XI3.XI3<6>.Y 0 0.101386f
c_73728 XI2.XI1.XI3.XI3<7>.NEN 0 0.0869923f
c_73746 XI2.XI1.XI3.XI3<6>.NEN 0 0.0876548f
c_73759 XI2.XI1.XI3.XI3<5>.X 0 0.0746321f
c_73773 XI2.XI1.XI3.XI3<4>.Y 0 0.100409f
c_73792 XI2.XI1.XI3.XI3<5>.NEN 0 0.086949f
c_73811 XI2.XI1.XI3.XI3<4>.NEN 0 0.0876263f
c_73826 XI2.XI1.XI3.XI3<10>.X 0 0.0750129f
c_73842 XI2.XI1.XI3.XI3<11>.Y 0 0.101556f
c_73856 XI2.XI1.XI3.XI3<11>.X 0 0.0743077f
c_73872 XI2.XI1.XI3.XI3<10>.Y 0 0.100781f
c_73891 XI2.XI1.XI3.XI3<11>.NEN 0 0.0871811f
c_73910 XI2.XI1.XI3.XI3<10>.NEN 0 0.0875662f
c_73924 XI2.XI1.XI3.XI3<9>.X 0 0.0749807f
c_73939 XI2.XI1.XI3.XI3<8>.Y 0 0.101368f
c_73957 XI2.XI1.XI3.XI3<9>.NEN 0 0.0871345f
c_73976 XI2.XI1.XI3.XI3<8>.NEN 0 0.0875624f
c_73992 XI2.XI1.XI3.XI3<14>.X 0 0.0718695f
c_74009 XI2.XI1.XI3.XI3<15>.Y 0 0.0998181f
c_74025 XI2.XI1.XI3.XI3<15>.X 0 0.072612f
c_74043 XI2.XI1.XI3.XI3<14>.Y 0 0.100032f
c_74061 XI2.XI1.XI3.XI3<15>.NEN 0 0.0876455f
c_74081 XI2.XI1.XI3.XI3<14>.NEN 0 0.0876004f
c_74095 XI2.XI1.XI3.XI3<13>.X 0 0.0732749f
c_74112 XI2.XI1.XI3.XI3<12>.Y 0 0.100921f
c_74132 XI2.XI1.XI3.XI3<13>.NEN 0 0.0869494f
c_74151 XI2.XI1.XI3.XI3<12>.NEN 0 0.0877192f
c_74166 XI2.XI1.XI4.XI3<4>.X 0 0.0749138f
c_74181 XI2.XI1.XI4.XI3<5>.Y 0 0.101787f
c_74196 XI2.XI1.XI4.XI3<8>.X 0 0.0741974f
c_74213 XI2.XI1.XI4.XI3<9>.Y 0 0.101197f
c_74230 XI2.XI1.XI4.XI3<12>.X 0 0.0725462f
c_74248 XI2.XI1.XI4.XI3<13>.Y 0 0.100511f
c_74262 XI2.XI1.XI4.XI3<2>.X 0 0.0747644f
c_74276 XI2.XI1.XI4.XI3<3>.Y 0 0.100903f
c_74289 XI2.XI1.XI4.XI3<3>.X 0 0.074512f
c_74303 XI2.XI1.XI4.XI3<2>.Y 0 0.100281f
c_74321 XI2.XI1.XI4.XI3<3>.NEN 0 0.0868931f
c_74339 XI2.XI1.XI4.XI3<2>.NEN 0 0.0876294f
c_74352 XI2.XI1.XI4.XI3<1>.X 0 0.0750365f
c_74365 XI2.XI1.XI4.XI3<0>.Y 0 0.102155f
c_74382 XI2.XI1.XI4.XI3<1>.NEN 0 0.0868938f
c_74398 XI2.XI1.XI4.XI3<0>.NEN 0 0.0881863f
c_74412 XI2.XI1.XI4.XI3<6>.X 0 0.0750161f
c_74428 XI2.XI1.XI4.XI3<7>.Y 0 0.100957f
c_74443 XI2.XI1.XI4.XI3<7>.X 0 0.0745502f
c_74459 XI2.XI1.XI4.XI3<6>.Y 0 0.101068f
c_74477 XI2.XI1.XI4.XI3<7>.NEN 0 0.0870956f
c_74496 XI2.XI1.XI4.XI3<6>.NEN 0 0.0875468f
c_74510 XI2.XI1.XI4.XI3<5>.X 0 0.0728477f
c_74525 XI2.XI1.XI4.XI3<4>.Y 0 0.100211f
c_74543 XI2.XI1.XI4.XI3<5>.NEN 0 0.0870708f
c_74562 XI2.XI1.XI4.XI3<4>.NEN 0 0.0875051f
c_74578 XI2.XI1.XI4.XI3<10>.X 0 0.0745514f
c_74595 XI2.XI1.XI4.XI3<11>.Y 0 0.101408f
c_74610 XI2.XI1.XI4.XI3<11>.X 0 0.0748205f
c_74627 XI2.XI1.XI4.XI3<10>.Y 0 0.100591f
c_74645 XI2.XI1.XI4.XI3<11>.NEN 0 0.0872244f
c_74664 XI2.XI1.XI4.XI3<10>.NEN 0 0.0875864f
c_74679 XI2.XI1.XI4.XI3<9>.X 0 0.0745491f
c_74695 XI2.XI1.XI4.XI3<8>.Y 0 0.101177f
c_74714 XI2.XI1.XI4.XI3<9>.NEN 0 0.0869342f
c_74733 XI2.XI1.XI4.XI3<8>.NEN 0 0.0875468f
c_74750 XI2.XI1.XI4.XI3<14>.X 0 0.0725454f
c_74768 XI2.XI1.XI4.XI3<15>.Y 0 0.100086f
c_74785 XI2.XI1.XI4.XI3<15>.X 0 0.0735599f
c_74804 XI2.XI1.XI4.XI3<14>.Y 0 0.100725f
c_74822 XI2.XI1.XI4.XI3<15>.NEN 0 0.0876464f
c_74842 XI2.XI1.XI4.XI3<14>.NEN 0 0.0875701f
c_74858 XI2.XI1.XI4.XI3<13>.X 0 0.0736412f
c_74876 XI2.XI1.XI4.XI3<12>.Y 0 0.101311f
c_74896 XI2.XI1.XI4.XI3<13>.NEN 0 0.086943f
c_74915 XI2.XI1.XI4.XI3<12>.NEN 0 0.0877414f
c_74930 XI2.XI1.XI6.XI3<0>.X 0 0.075315f
c_74943 XI2.XI1.XI6.XI3<1>.Y 0 0.100947f
c_74957 XI2.XI1.XI6.XI3<4>.X 0 0.0747698f
c_74972 XI2.XI1.XI6.XI3<5>.Y 0 0.10152f
c_74987 XI2.XI1.XI6.XI3<8>.X 0 0.0748546f
c_75003 XI2.XI1.XI6.XI3<9>.Y 0 0.101356f
c_75020 XI2.XI1.XI6.XI3<12>.X 0 0.07287f
c_75038 XI2.XI1.XI6.XI3<13>.Y 0 0.100511f
c_75052 XI2.XI1.XI6.XI3<2>.X 0 0.0750422f
c_75066 XI2.XI1.XI6.XI3<3>.Y 0 0.100901f
c_75079 XI2.XI1.XI6.XI3<3>.X 0 0.0745673f
c_75093 XI2.XI1.XI6.XI3<2>.Y 0 0.100306f
c_75111 XI2.XI1.XI6.XI3<3>.NEN 0 0.0868931f
c_75129 XI2.XI1.XI6.XI3<2>.NEN 0 0.0876294f
c_75142 XI2.XI1.XI6.XI3<1>.X 0 0.0750372f
c_75155 XI2.XI1.XI6.XI3<0>.Y 0 0.102164f
c_75172 XI2.XI1.XI6.XI3<1>.NEN 0 0.0868938f
c_75188 XI2.XI1.XI6.XI3<0>.NEN 0 0.0882254f
c_75202 XI2.XI1.XI6.XI3<6>.X 0 0.0752697f
c_75218 XI2.XI1.XI6.XI3<7>.Y 0 0.101434f
c_75233 XI2.XI1.XI6.XI3<7>.X 0 0.0749457f
c_75248 XI2.XI1.XI6.XI3<6>.Y 0 0.101231f
c_75266 XI2.XI1.XI6.XI3<7>.NEN 0 0.0871095f
c_75285 XI2.XI1.XI6.XI3<6>.NEN 0 0.0875468f
c_75299 XI2.XI1.XI6.XI3<5>.X 0 0.0749434f
c_75314 XI2.XI1.XI6.XI3<4>.Y 0 0.100212f
c_75332 XI2.XI1.XI6.XI3<5>.NEN 0 0.087056f
c_75351 XI2.XI1.XI6.XI3<4>.NEN 0 0.0874208f
c_75367 XI2.XI1.XI6.XI3<10>.X 0 0.0748381f
c_75384 XI2.XI1.XI6.XI3<11>.Y 0 0.100952f
c_75399 XI2.XI1.XI6.XI3<11>.X 0 0.0748016f
c_75416 XI2.XI1.XI6.XI3<10>.Y 0 0.10059f
c_75435 XI2.XI1.XI6.XI3<11>.NEN 0 0.0871728f
c_75454 XI2.XI1.XI6.XI3<10>.NEN 0 0.0875864f
c_75469 XI2.XI1.XI6.XI3<9>.X 0 0.0745574f
c_75485 XI2.XI1.XI6.XI3<8>.Y 0 0.101236f
c_75504 XI2.XI1.XI6.XI3<9>.NEN 0 0.0869342f
c_75523 XI2.XI1.XI6.XI3<8>.NEN 0 0.087563f
c_75540 XI2.XI1.XI6.XI3<14>.X 0 0.0723887f
c_75558 XI2.XI1.XI6.XI3<15>.Y 0 0.100086f
c_75575 XI2.XI1.XI6.XI3<15>.X 0 0.0735654f
c_75594 XI2.XI1.XI6.XI3<14>.Y 0 0.100565f
c_75612 XI2.XI1.XI6.XI3<15>.NEN 0 0.0876766f
c_75632 XI2.XI1.XI6.XI3<14>.NEN 0 0.0875701f
c_75648 XI2.XI1.XI6.XI3<13>.X 0 0.0736484f
c_75666 XI2.XI1.XI6.XI3<12>.Y 0 0.101311f
c_75686 XI2.XI1.XI6.XI3<13>.NEN 0 0.086943f
c_75705 XI2.XI1.XI6.XI3<12>.NEN 0 0.0877414f
c_75719 XI2.XI1.XI5.XI3<4>.X 0 0.0747648f
c_75734 XI2.XI1.XI5.XI3<5>.Y 0 0.10152f
c_75749 XI2.XI1.XI5.XI3<8>.X 0 0.0748546f
c_75765 XI2.XI1.XI5.XI3<9>.Y 0 0.101356f
c_75781 XI2.XI1.XI5.XI3<12>.X 0 0.0728928f
c_75799 XI2.XI1.XI5.XI3<13>.Y 0 0.100511f
c_75813 XI2.XI1.XI5.XI3<2>.X 0 0.0785812f
c_75827 XI2.XI1.XI5.XI3<3>.Y 0 0.101098f
c_75840 XI2.XI1.XI5.XI3<3>.X 0 0.0756793f
c_75854 XI2.XI1.XI5.XI3<2>.Y 0 0.102053f
c_75872 XI2.XI1.XI5.XI3<3>.NEN 0 0.0868931f
c_75890 XI2.XI1.XI5.XI3<2>.NEN 0 0.0876223f
c_75903 XI2.XI1.XI5.XI3<1>.X 0 0.0749568f
c_75917 XI2.XI1.XI5.XI3<0>.Y 0 0.101991f
c_75934 XI2.XI1.XI5.XI3<1>.NEN 0 0.0868938f
c_75951 XI2.XI1.XI5.XI3<0>.NEN 0 0.0881404f
c_75965 XI2.XI1.XI5.XI3<6>.X 0 0.0752697f
c_75981 XI2.XI1.XI5.XI3<7>.Y 0 0.101401f
c_75996 XI2.XI1.XI5.XI3<7>.X 0 0.0749457f
c_76011 XI2.XI1.XI5.XI3<6>.Y 0 0.101231f
c_76029 XI2.XI1.XI5.XI3<7>.NEN 0 0.0871095f
c_76048 XI2.XI1.XI5.XI3<6>.NEN 0 0.0875468f
c_76062 XI2.XI1.XI5.XI3<5>.X 0 0.0749434f
c_76077 XI2.XI1.XI5.XI3<4>.Y 0 0.100214f
c_76095 XI2.XI1.XI5.XI3<5>.NEN 0 0.087056f
c_76113 XI2.XI1.XI5.XI3<4>.NEN 0 0.0875193f
c_76129 XI2.XI1.XI5.XI3<10>.X 0 0.0748381f
c_76146 XI2.XI1.XI5.XI3<11>.Y 0 0.101303f
c_76161 XI2.XI1.XI5.XI3<11>.X 0 0.0748016f
c_76178 XI2.XI1.XI5.XI3<10>.Y 0 0.100589f
c_76197 XI2.XI1.XI5.XI3<11>.NEN 0 0.0871719f
c_76216 XI2.XI1.XI5.XI3<10>.NEN 0 0.0875864f
c_76231 XI2.XI1.XI5.XI3<9>.X 0 0.0745574f
c_76247 XI2.XI1.XI5.XI3<8>.Y 0 0.101236f
c_76266 XI2.XI1.XI5.XI3<9>.NEN 0 0.0869342f
c_76285 XI2.XI1.XI5.XI3<8>.NEN 0 0.0875767f
c_76302 XI2.XI1.XI5.XI3<14>.X 0 0.0723887f
c_76320 XI2.XI1.XI5.XI3<15>.Y 0 0.100004f
c_76337 XI2.XI1.XI5.XI3<15>.X 0 0.073566f
c_76355 XI2.XI1.XI5.XI3<14>.Y 0 0.100728f
c_76373 XI2.XI1.XI5.XI3<15>.NEN 0 0.0876716f
c_76393 XI2.XI1.XI5.XI3<14>.NEN 0 0.0875701f
c_76409 XI2.XI1.XI5.XI3<13>.X 0 0.0736484f
c_76427 XI2.XI1.XI5.XI3<12>.Y 0 0.101311f
c_76447 XI2.XI1.XI5.XI3<13>.NEN 0 0.086947f
c_76466 XI2.XI1.XI5.XI3<12>.NEN 0 0.0877414f
c_76481 XI2.XI1.XI10.XI3<0>.X 0 0.0753166f
c_76494 XI2.XI1.XI10.XI3<1>.Y 0 0.100839f
c_76508 XI2.XI1.XI10.XI3<4>.X 0 0.0747648f
c_76523 XI2.XI1.XI10.XI3<5>.Y 0 0.101511f
c_76538 XI2.XI1.XI10.XI3<8>.X 0 0.0748546f
c_76554 XI2.XI1.XI10.XI3<9>.Y 0 0.10305f
c_76570 XI2.XI1.XI10.XI3<12>.X 0 0.0728928f
c_76588 XI2.XI1.XI10.XI3<13>.Y 0 0.100511f
c_76602 XI2.XI1.XI10.XI3<2>.X 0 0.0785692f
c_76616 XI2.XI1.XI10.XI3<3>.Y 0 0.100814f
c_76629 XI2.XI1.XI10.XI3<3>.X 0 0.0757948f
c_76643 XI2.XI1.XI10.XI3<2>.Y 0 0.102053f
c_76661 XI2.XI1.XI10.XI3<3>.NEN 0 0.0868951f
c_76679 XI2.XI1.XI10.XI3<2>.NEN 0 0.0875051f
c_76691 XI2.XI1.XI10.XI3<1>.X 0 0.0754703f
c_76705 XI2.XI1.XI10.XI3<0>.Y 0 0.102032f
c_76722 XI2.XI1.XI10.XI3<1>.NEN 0 0.0868938f
c_76739 XI2.XI1.XI10.XI3<0>.NEN 0 0.0882325f
c_76753 XI2.XI1.XI10.XI3<6>.X 0 0.0753324f
c_76769 XI2.XI1.XI10.XI3<7>.Y 0 0.101317f
c_76784 XI2.XI1.XI10.XI3<7>.X 0 0.0749457f
c_76799 XI2.XI1.XI10.XI3<6>.Y 0 0.10126f
c_76817 XI2.XI1.XI10.XI3<7>.NEN 0 0.0871095f
c_76836 XI2.XI1.XI10.XI3<6>.NEN 0 0.0875468f
c_76850 XI2.XI1.XI10.XI3<5>.X 0 0.07494f
c_76865 XI2.XI1.XI10.XI3<4>.Y 0 0.100058f
c_76883 XI2.XI1.XI10.XI3<5>.NEN 0 0.087056f
c_76901 XI2.XI1.XI10.XI3<4>.NEN 0 0.0875193f
c_76917 XI2.XI1.XI10.XI3<10>.X 0 0.0748381f
c_76934 XI2.XI1.XI10.XI3<11>.Y 0 0.101464f
c_76949 XI2.XI1.XI10.XI3<11>.X 0 0.0748016f
c_76966 XI2.XI1.XI10.XI3<10>.Y 0 0.100589f
c_76985 XI2.XI1.XI10.XI3<11>.NEN 0 0.0871714f
c_77004 XI2.XI1.XI10.XI3<10>.NEN 0 0.0875792f
c_77019 XI2.XI1.XI10.XI3<9>.X 0 0.0736655f
c_77035 XI2.XI1.XI10.XI3<8>.Y 0 0.101236f
c_77054 XI2.XI1.XI10.XI3<9>.NEN 0 0.0869529f
c_77073 XI2.XI1.XI10.XI3<8>.NEN 0 0.0875767f
c_77090 XI2.XI1.XI10.XI3<14>.X 0 0.0723887f
c_77108 XI2.XI1.XI10.XI3<15>.Y 0 0.0999863f
c_77125 XI2.XI1.XI10.XI3<15>.X 0 0.0735666f
c_77143 XI2.XI1.XI10.XI3<14>.Y 0 0.100728f
c_77161 XI2.XI1.XI10.XI3<15>.NEN 0 0.0876091f
c_77181 XI2.XI1.XI10.XI3<14>.NEN 0 0.0875701f
c_77198 XI2.XI1.XI10.XI3<13>.X 0 0.073538f
c_77216 XI2.XI1.XI10.XI3<12>.Y 0 0.101308f
c_77236 XI2.XI1.XI10.XI3<13>.NEN 0 0.086947f
c_77255 XI2.XI1.XI10.XI3<12>.NEN 0 0.087729f
c_77269 XI2.XI1.XI9.XI3<4>.X 0 0.0752609f
c_77284 XI2.XI1.XI9.XI3<5>.Y 0 0.101477f
c_77299 XI2.XI1.XI9.XI3<8>.X 0 0.0748546f
c_77315 XI2.XI1.XI9.XI3<9>.Y 0 0.103525f
c_77331 XI2.XI1.XI9.XI3<12>.X 0 0.0728928f
c_77349 XI2.XI1.XI9.XI3<13>.Y 0 0.100502f
c_77362 XI2.XI1.XI9.XI3<2>.X 0 0.0784206f
c_77376 XI2.XI1.XI9.XI3<3>.Y 0 0.100812f
c_77389 XI2.XI1.XI9.XI3<3>.X 0 0.0758441f
c_77403 XI2.XI1.XI9.XI3<2>.Y 0 0.102053f
c_77421 XI2.XI1.XI9.XI3<3>.NEN 0 0.0868992f
c_77439 XI2.XI1.XI9.XI3<2>.NEN 0 0.0874208f
c_77451 XI2.XI1.XI9.XI3<1>.X 0 0.0751195f
c_77465 XI2.XI1.XI9.XI3<0>.Y 0 0.102112f
c_77482 XI2.XI1.XI9.XI3<1>.NEN 0 0.0868938f
c_77499 XI2.XI1.XI9.XI3<0>.NEN 0 0.0881863f
c_77514 XI2.XI1.XI9.XI3<6>.X 0 0.0748347f
c_77529 XI2.XI1.XI9.XI3<7>.Y 0 0.101476f
c_77544 XI2.XI1.XI9.XI3<7>.X 0 0.0749491f
c_77559 XI2.XI1.XI9.XI3<6>.Y 0 0.101266f
c_77577 XI2.XI1.XI9.XI3<7>.NEN 0 0.0869906f
c_77596 XI2.XI1.XI9.XI3<6>.NEN 0 0.0875468f
c_77610 XI2.XI1.XI9.XI3<5>.X 0 0.07494f
c_77624 XI2.XI1.XI9.XI3<4>.Y 0 0.100218f
c_77642 XI2.XI1.XI9.XI3<5>.NEN 0 0.087001f
c_77660 XI2.XI1.XI9.XI3<4>.NEN 0 0.0875193f
c_77676 XI2.XI1.XI9.XI3<10>.X 0 0.0748381f
c_77693 XI2.XI1.XI9.XI3<11>.Y 0 0.101462f
c_77708 XI2.XI1.XI9.XI3<11>.X 0 0.0748016f
c_77725 XI2.XI1.XI9.XI3<10>.Y 0 0.10059f
c_77744 XI2.XI1.XI9.XI3<11>.NEN 0 0.0871733f
c_77763 XI2.XI1.XI9.XI3<10>.NEN 0 0.0875721f
c_77777 XI2.XI1.XI9.XI3<9>.X 0 0.0737546f
c_77793 XI2.XI1.XI9.XI3<8>.Y 0 0.101235f
c_77812 XI2.XI1.XI9.XI3<9>.NEN 0 0.0869859f
c_77831 XI2.XI1.XI9.XI3<8>.NEN 0 0.0875767f
c_77848 XI2.XI1.XI9.XI3<14>.X 0 0.0723887f
c_77866 XI2.XI1.XI9.XI3<15>.Y 0 0.0999109f
c_77883 XI2.XI1.XI9.XI3<15>.X 0 0.0735664f
c_77901 XI2.XI1.XI9.XI3<14>.Y 0 0.100728f
c_77919 XI2.XI1.XI9.XI3<15>.NEN 0 0.0875356f
c_77939 XI2.XI1.XI9.XI3<14>.NEN 0 0.0875701f
c_77955 XI2.XI1.XI9.XI3<13>.X 0 0.0738007f
c_77973 XI2.XI1.XI9.XI3<12>.Y 0 0.101148f
c_77993 XI2.XI1.XI9.XI3<13>.NEN 0 0.086947f
c_78012 XI2.XI1.XI9.XI3<12>.NEN 0 0.087729f
c_78027 XI2.XI1.XI7.XI3<0>.X 0 0.0753064f
c_78041 XI2.XI1.XI7.XI3<1>.Y 0 0.100762f
c_78055 XI2.XI1.XI7.XI3<4>.X 0 0.0752787f
c_78070 XI2.XI1.XI7.XI3<5>.Y 0 0.101353f
c_78085 XI2.XI1.XI7.XI3<8>.X 0 0.0748543f
c_78101 XI2.XI1.XI7.XI3<9>.Y 0 0.101959f
c_78117 XI2.XI1.XI7.XI3<12>.X 0 0.0728928f
c_78135 XI2.XI1.XI7.XI3<13>.Y 0 0.100469f
c_78148 XI2.XI1.XI7.XI3<2>.X 0 0.0784206f
c_78162 XI2.XI1.XI7.XI3<3>.Y 0 0.100813f
c_78176 XI2.XI1.XI7.XI3<3>.X 0 0.075737f
c_78190 XI2.XI1.XI7.XI3<2>.Y 0 0.102049f
c_78208 XI2.XI1.XI7.XI3<3>.NEN 0 0.0868992f
c_78225 XI2.XI1.XI7.XI3<2>.NEN 0 0.0875193f
c_78237 XI2.XI1.XI7.XI3<1>.X 0 0.0750456f
c_78251 XI2.XI1.XI7.XI3<0>.Y 0 0.102147f
c_78268 XI2.XI1.XI7.XI3<1>.NEN 0 0.0868938f
c_78285 XI2.XI1.XI7.XI3<0>.NEN 0 0.0881863f
c_78300 XI2.XI1.XI7.XI3<6>.X 0 0.0748347f
c_78315 XI2.XI1.XI7.XI3<7>.Y 0 0.101475f
c_78330 XI2.XI1.XI7.XI3<7>.X 0 0.0749491f
c_78345 XI2.XI1.XI7.XI3<6>.Y 0 0.101266f
c_78363 XI2.XI1.XI7.XI3<7>.NEN 0 0.0869906f
c_78382 XI2.XI1.XI7.XI3<6>.NEN 0 0.0875468f
c_78396 XI2.XI1.XI7.XI3<5>.X 0 0.0749998f
c_78410 XI2.XI1.XI7.XI3<4>.Y 0 0.100218f
c_78428 XI2.XI1.XI7.XI3<5>.NEN 0 0.0870009f
c_78446 XI2.XI1.XI7.XI3<4>.NEN 0 0.0875193f
c_78462 XI2.XI1.XI7.XI3<10>.X 0 0.0748233f
c_78479 XI2.XI1.XI7.XI3<11>.Y 0 0.101461f
c_78494 XI2.XI1.XI7.XI3<11>.X 0 0.0748016f
c_78511 XI2.XI1.XI7.XI3<10>.Y 0 0.10059f
c_78530 XI2.XI1.XI7.XI3<11>.NEN 0 0.0871905f
c_78549 XI2.XI1.XI7.XI3<10>.NEN 0 0.0874878f
c_78563 XI2.XI1.XI7.XI3<9>.X 0 0.0743231f
c_78579 XI2.XI1.XI7.XI3<8>.Y 0 0.101235f
c_78598 XI2.XI1.XI7.XI3<9>.NEN 0 0.0869859f
c_78617 XI2.XI1.XI7.XI3<8>.NEN 0 0.0875767f
c_78635 XI2.XI1.XI7.XI3<14>.X 0 0.0723887f
c_78652 XI2.XI1.XI7.XI3<15>.Y 0 0.100091f
c_78669 XI2.XI1.XI7.XI3<15>.X 0 0.0735657f
c_78687 XI2.XI1.XI7.XI3<14>.Y 0 0.100728f
c_78704 XI2.XI1.XI7.XI3<15>.NEN 0 0.0876798f
c_78724 XI2.XI1.XI7.XI3<14>.NEN 0 0.0875701f
c_78740 XI2.XI1.XI7.XI3<13>.X 0 0.0738007f
c_78757 XI2.XI1.XI7.XI3<12>.Y 0 0.101311f
c_78777 XI2.XI1.XI7.XI3<13>.NEN 0 0.086947f
c_78796 XI2.XI1.XI7.XI3<12>.NEN 0 0.087729f
c_78810 XI2.XI1.XI8.XI3<4>.X 0 0.0752991f
c_78825 XI2.XI1.XI8.XI3<5>.Y 0 0.101269f
c_78840 XI2.XI1.XI8.XI3<8>.X 0 0.0748437f
c_78856 XI2.XI1.XI8.XI3<9>.Y 0 0.101963f
c_78872 XI2.XI1.XI8.XI3<12>.X 0 0.0728928f
c_78890 XI2.XI1.XI8.XI3<13>.Y 0 0.100437f
c_78903 XI2.XI1.XI8.XI3<2>.X 0 0.0784206f
c_78917 XI2.XI1.XI8.XI3<3>.Y 0 0.100804f
c_78930 XI2.XI1.XI8.XI3<3>.X 0 0.0769124f
c_78944 XI2.XI1.XI8.XI3<2>.Y 0 0.101895f
c_78962 XI2.XI1.XI8.XI3<3>.NEN 0 0.0868992f
c_78979 XI2.XI1.XI8.XI3<2>.NEN 0 0.0875193f
c_78991 XI2.XI1.XI8.XI3<1>.X 0 0.0750456f
c_79005 XI2.XI1.XI8.XI3<0>.Y 0 0.102198f
c_79022 XI2.XI1.XI8.XI3<1>.NEN 0 0.0868938f
c_79039 XI2.XI1.XI8.XI3<0>.NEN 0 0.0882353f
c_79054 XI2.XI1.XI8.XI3<6>.X 0 0.0748347f
c_79069 XI2.XI1.XI8.XI3<7>.Y 0 0.101475f
c_79084 XI2.XI1.XI8.XI3<7>.X 0 0.07486f
c_79099 XI2.XI1.XI8.XI3<6>.Y 0 0.101266f
c_79117 XI2.XI1.XI8.XI3<7>.NEN 0 0.0869906f
c_79136 XI2.XI1.XI8.XI3<6>.NEN 0 0.0875468f
c_79150 XI2.XI1.XI8.XI3<5>.X 0 0.0749998f
c_79164 XI2.XI1.XI8.XI3<4>.Y 0 0.100243f
c_79182 XI2.XI1.XI8.XI3<5>.NEN 0 0.0870009f
c_79200 XI2.XI1.XI8.XI3<4>.NEN 0 0.0875193f
c_79216 XI2.XI1.XI8.XI3<10>.X 0 0.0748233f
c_79233 XI2.XI1.XI8.XI3<11>.Y 0 0.101462f
c_79248 XI2.XI1.XI8.XI3<11>.X 0 0.0748016f
c_79265 XI2.XI1.XI8.XI3<10>.Y 0 0.100586f
c_79284 XI2.XI1.XI8.XI3<11>.NEN 0 0.0871762f
c_79302 XI2.XI1.XI8.XI3<10>.NEN 0 0.0875864f
c_79316 XI2.XI1.XI8.XI3<9>.X 0 0.0750082f
c_79332 XI2.XI1.XI8.XI3<8>.Y 0 0.101235f
c_79351 XI2.XI1.XI8.XI3<9>.NEN 0 0.0869859f
c_79370 XI2.XI1.XI8.XI3<8>.NEN 0 0.0875767f
c_79388 XI2.XI1.XI8.XI3<14>.X 0 0.0723887f
c_79405 XI2.XI1.XI8.XI3<15>.Y 0 0.100119f
c_79422 XI2.XI1.XI8.XI3<15>.X 0 0.0735656f
c_79440 XI2.XI1.XI8.XI3<14>.Y 0 0.100728f
c_79457 XI2.XI1.XI8.XI3<15>.NEN 0 0.0876589f
c_79477 XI2.XI1.XI8.XI3<14>.NEN 0 0.0875701f
c_79493 XI2.XI1.XI8.XI3<13>.X 0 0.0738007f
c_79510 XI2.XI1.XI8.XI3<12>.Y 0 0.101311f
c_79530 XI2.XI1.XI8.XI3<13>.NEN 0 0.086947f
c_79549 XI2.XI1.XI8.XI3<12>.NEN 0 0.087729f
c_79563 XI2.XI1.XI11.XI3<0>.X 0 0.0753144f
c_79577 XI2.XI1.XI11.XI3<1>.Y 0 0.100947f
c_79591 XI2.XI1.XI11.XI3<4>.X 0 0.0752871f
c_79605 XI2.XI1.XI11.XI3<5>.Y 0 0.10152f
c_79620 XI2.XI1.XI11.XI3<8>.X 0 0.0748317f
c_79636 XI2.XI1.XI11.XI3<9>.Y 0 0.101963f
c_79652 XI2.XI1.XI11.XI3<12>.X 0 0.0728928f
c_79670 XI2.XI1.XI11.XI3<13>.Y 0 0.10035f
c_79683 XI2.XI1.XI11.XI3<2>.X 0 0.0784206f
c_79697 XI2.XI1.XI11.XI3<3>.Y 0 0.102987f
c_79710 XI2.XI1.XI11.XI3<3>.X 0 0.076201f
c_79723 XI2.XI1.XI11.XI3<2>.Y 0 0.102053f
c_79741 XI2.XI1.XI11.XI3<3>.NEN 0 0.0868992f
c_79758 XI2.XI1.XI11.XI3<2>.NEN 0 0.0875193f
c_79770 XI2.XI1.XI11.XI3<1>.X 0 0.0750456f
c_79784 XI2.XI1.XI11.XI3<0>.Y 0 0.10221f
c_79802 XI2.XI1.XI11.XI3<1>.NEN 0 0.0867791f
c_79820 XI2.XI1.XI11.XI3<0>.NEN 0 0.0879949f
c_79835 XI2.XI1.XI11.XI3<6>.X 0 0.0748347f
c_79850 XI2.XI1.XI11.XI3<7>.Y 0 0.101475f
c_79864 XI2.XI1.XI11.XI3<7>.X 0 0.0749491f
c_79879 XI2.XI1.XI11.XI3<6>.Y 0 0.101266f
c_79897 XI2.XI1.XI11.XI3<7>.NEN 0 0.0870011f
c_79916 XI2.XI1.XI11.XI3<6>.NEN 0 0.0875468f
c_79930 XI2.XI1.XI11.XI3<5>.X 0 0.0749362f
c_79944 XI2.XI1.XI11.XI3<4>.Y 0 0.10028f
c_79962 XI2.XI1.XI11.XI3<5>.NEN 0 0.0868938f
c_79980 XI2.XI1.XI11.XI3<4>.NEN 0 0.0875193f
c_79996 XI2.XI1.XI11.XI3<10>.X 0 0.0748233f
c_80013 XI2.XI1.XI11.XI3<11>.Y 0 0.101909f
c_80028 XI2.XI1.XI11.XI3<11>.X 0 0.0748016f
c_80045 XI2.XI1.XI11.XI3<10>.Y 0 0.100425f
c_80064 XI2.XI1.XI11.XI3<11>.NEN 0 0.0871757f
c_80082 XI2.XI1.XI11.XI3<10>.NEN 0 0.0875864f
c_80096 XI2.XI1.XI11.XI3<9>.X 0 0.0750237f
c_80112 XI2.XI1.XI11.XI3<8>.Y 0 0.101235f
c_80131 XI2.XI1.XI11.XI3<9>.NEN 0 0.0869859f
c_80150 XI2.XI1.XI11.XI3<8>.NEN 0 0.0875767f
c_80168 XI2.XI1.XI11.XI3<14>.X 0 0.0723887f
c_80185 XI2.XI1.XI11.XI3<15>.Y 0 0.100048f
c_80202 XI2.XI1.XI11.XI3<15>.X 0 0.0735663f
c_80221 XI2.XI1.XI11.XI3<14>.Y 0 0.100541f
c_80238 XI2.XI1.XI11.XI3<15>.NEN 0 0.0877016f
c_80258 XI2.XI1.XI11.XI3<14>.NEN 0 0.0875826f
c_80274 XI2.XI1.XI11.XI3<13>.X 0 0.0738007f
c_80291 XI2.XI1.XI11.XI3<12>.Y 0 0.101311f
c_80311 XI2.XI1.XI11.XI3<13>.NEN 0 0.0869449f
c_80330 XI2.XI1.XI11.XI3<12>.NEN 0 0.087729f
c_80344 XI2.XI1.XI12.XI3<4>.X 0 0.0752871f
c_80358 XI2.XI1.XI12.XI3<5>.Y 0 0.101519f
c_80372 XI2.XI1.XI12.XI3<8>.X 0 0.0748546f
c_80388 XI2.XI1.XI12.XI3<9>.Y 0 0.101963f
c_80405 XI2.XI1.XI12.XI3<12>.X 0 0.0728928f
c_80422 XI2.XI1.XI12.XI3<13>.Y 0 0.100511f
c_80435 XI2.XI1.XI12.XI3<2>.X 0 0.0784256f
c_80449 XI2.XI1.XI12.XI3<3>.Y 0 0.102955f
c_80462 XI2.XI1.XI12.XI3<3>.X 0 0.0765056f
c_80475 XI2.XI1.XI12.XI3<2>.Y 0 0.10246f
c_80493 XI2.XI1.XI12.XI3<3>.NEN 0 0.0868992f
c_80510 XI2.XI1.XI12.XI3<2>.NEN 0 0.0875193f
c_80523 XI2.XI1.XI12.XI3<1>.X 0 0.0749419f
c_80537 XI2.XI1.XI12.XI3<0>.Y 0 0.102175f
c_80555 XI2.XI1.XI12.XI3<1>.NEN 0 0.0868526f
c_80572 XI2.XI1.XI12.XI3<0>.NEN 0 0.0881263f
c_80587 XI2.XI1.XI12.XI3<6>.X 0 0.0748347f
c_80602 XI2.XI1.XI12.XI3<7>.Y 0 0.101552f
c_80616 XI2.XI1.XI12.XI3<7>.X 0 0.0749491f
c_80631 XI2.XI1.XI12.XI3<6>.Y 0 0.101265f
c_80649 XI2.XI1.XI12.XI3<7>.NEN 0 0.0870022f
c_80668 XI2.XI1.XI12.XI3<6>.NEN 0 0.0875468f
c_80682 XI2.XI1.XI12.XI3<5>.X 0 0.0749362f
c_80696 XI2.XI1.XI12.XI3<4>.Y 0 0.10028f
c_80714 XI2.XI1.XI12.XI3<5>.NEN 0 0.0868938f
c_80732 XI2.XI1.XI12.XI3<4>.NEN 0 0.0875193f
c_80748 XI2.XI1.XI12.XI3<10>.X 0 0.0748233f
c_80765 XI2.XI1.XI12.XI3<11>.Y 0 0.101876f
c_80780 XI2.XI1.XI12.XI3<11>.X 0 0.0748016f
c_80796 XI2.XI1.XI12.XI3<10>.Y 0 0.100588f
c_80815 XI2.XI1.XI12.XI3<11>.NEN 0 0.0871742f
c_80833 XI2.XI1.XI12.XI3<10>.NEN 0 0.0875864f
c_80847 XI2.XI1.XI12.XI3<9>.X 0 0.0754565f
c_80863 XI2.XI1.XI12.XI3<8>.Y 0 0.101235f
c_80882 XI2.XI1.XI12.XI3<9>.NEN 0 0.0869866f
c_80901 XI2.XI1.XI12.XI3<8>.NEN 0 0.0875767f
c_80919 XI2.XI1.XI12.XI3<14>.X 0 0.0723887f
c_80936 XI2.XI1.XI12.XI3<15>.Y 0 0.100064f
c_80953 XI2.XI1.XI12.XI3<15>.X 0 0.0735248f
c_80972 XI2.XI1.XI12.XI3<14>.Y 0 0.100617f
c_80989 XI2.XI1.XI12.XI3<15>.NEN 0 0.0876148f
c_81009 XI2.XI1.XI12.XI3<14>.NEN 0 0.0875826f
c_81025 XI2.XI1.XI12.XI3<13>.X 0 0.0738007f
c_81042 XI2.XI1.XI12.XI3<12>.Y 0 0.101311f
c_81062 XI2.XI1.XI12.XI3<13>.NEN 0 0.0869356f
c_81081 XI2.XI1.XI12.XI3<12>.NEN 0 0.087729f
c_81095 XI2.XI1.XI14.XI3<0>.X 0 0.0753192f
c_81109 XI2.XI1.XI14.XI3<1>.Y 0 0.100947f
c_81123 XI2.XI1.XI14.XI3<4>.X 0 0.0752871f
c_81137 XI2.XI1.XI14.XI3<5>.Y 0 0.10152f
c_81151 XI2.XI1.XI14.XI3<8>.X 0 0.0748546f
c_81167 XI2.XI1.XI14.XI3<9>.Y 0 0.101963f
c_81184 XI2.XI1.XI14.XI3<12>.X 0 0.0728928f
c_81201 XI2.XI1.XI14.XI3<13>.Y 0 0.100511f
c_81214 XI2.XI1.XI14.XI3<2>.X 0 0.0747644f
c_81228 XI2.XI1.XI14.XI3<3>.Y 0 0.102872f
c_81242 XI2.XI1.XI14.XI3<3>.X 0 0.07528f
c_81255 XI2.XI1.XI14.XI3<2>.Y 0 0.100281f
c_81273 XI2.XI1.XI14.XI3<3>.NEN 0 0.0868257f
c_81290 XI2.XI1.XI14.XI3<2>.NEN 0 0.0875193f
c_81303 XI2.XI1.XI14.XI3<1>.X 0 0.0750284f
c_81317 XI2.XI1.XI14.XI3<0>.Y 0 0.102034f
c_81335 XI2.XI1.XI14.XI3<1>.NEN 0 0.086883f
c_81352 XI2.XI1.XI14.XI3<0>.NEN 0 0.0880698f
c_81367 XI2.XI1.XI14.XI3<6>.X 0 0.0748238f
c_81382 XI2.XI1.XI14.XI3<7>.Y 0 0.10158f
c_81396 XI2.XI1.XI14.XI3<7>.X 0 0.0749491f
c_81411 XI2.XI1.XI14.XI3<6>.Y 0 0.101266f
c_81429 XI2.XI1.XI14.XI3<7>.NEN 0 0.0870033f
c_81448 XI2.XI1.XI14.XI3<6>.NEN 0 0.0875397f
c_81462 XI2.XI1.XI14.XI3<5>.X 0 0.0748471f
c_81477 XI2.XI1.XI14.XI3<4>.Y 0 0.100097f
c_81495 XI2.XI1.XI14.XI3<5>.NEN 0 0.0868938f
c_81513 XI2.XI1.XI14.XI3<4>.NEN 0 0.0875193f
c_81529 XI2.XI1.XI14.XI3<10>.X 0 0.0748233f
c_81546 XI2.XI1.XI14.XI3<11>.Y 0 0.101387f
c_81561 XI2.XI1.XI14.XI3<11>.X 0 0.0748016f
c_81577 XI2.XI1.XI14.XI3<10>.Y 0 0.100588f
c_81596 XI2.XI1.XI14.XI3<11>.NEN 0 0.0871723f
c_81614 XI2.XI1.XI14.XI3<10>.NEN 0 0.0875864f
c_81628 XI2.XI1.XI14.XI3<9>.X 0 0.0754565f
c_81644 XI2.XI1.XI14.XI3<8>.Y 0 0.101231f
c_81663 XI2.XI1.XI14.XI3<9>.NEN 0 0.0869866f
c_81682 XI2.XI1.XI14.XI3<8>.NEN 0 0.0875468f
c_81700 XI2.XI1.XI14.XI3<14>.X 0 0.0723887f
c_81717 XI2.XI1.XI14.XI3<15>.Y 0 0.100088f
c_81734 XI2.XI1.XI14.XI3<15>.X 0 0.0735244f
c_81753 XI2.XI1.XI14.XI3<14>.Y 0 0.100677f
c_81770 XI2.XI1.XI14.XI3<15>.NEN 0 0.0876091f
c_81790 XI2.XI1.XI14.XI3<14>.NEN 0 0.0875826f
c_81806 XI2.XI1.XI14.XI3<13>.X 0 0.0738007f
c_81823 XI2.XI1.XI14.XI3<12>.Y 0 0.101311f
c_81843 XI2.XI1.XI14.XI3<13>.NEN 0 0.0869356f
c_81862 XI2.XI1.XI14.XI3<12>.NEN 0 0.087729f
c_81876 XI2.XI1.XI13.XI3<4>.X 0 0.0752871f
c_81890 XI2.XI1.XI13.XI3<5>.Y 0 0.10152f
c_81904 XI2.XI1.XI13.XI3<8>.X 0 0.0748546f
c_81920 XI2.XI1.XI13.XI3<9>.Y 0 0.101955f
c_81937 XI2.XI1.XI13.XI3<12>.X 0 0.0728928f
c_81954 XI2.XI1.XI13.XI3<13>.Y 0 0.100511f
c_81968 XI2.XI1.XI13.XI3<2>.X 0 0.0784206f
c_81981 XI2.XI1.XI13.XI3<3>.Y 0 0.103171f
c_81994 XI2.XI1.XI13.XI3<3>.X 0 0.0780287f
c_82007 XI2.XI1.XI13.XI3<2>.Y 0 0.102053f
c_82024 XI2.XI1.XI13.XI3<3>.NEN 0 0.0868992f
c_82041 XI2.XI1.XI13.XI3<2>.NEN 0 0.0875193f
c_82054 XI2.XI1.XI13.XI3<1>.X 0 0.0750456f
c_82067 XI2.XI1.XI13.XI3<0>.Y 0 0.102194f
c_82085 XI2.XI1.XI13.XI3<1>.NEN 0 0.0868938f
c_82102 XI2.XI1.XI13.XI3<0>.NEN 0 0.0880683f
c_82117 XI2.XI1.XI13.XI3<6>.X 0 0.0748117f
c_82132 XI2.XI1.XI13.XI3<7>.Y 0 0.101574f
c_82146 XI2.XI1.XI13.XI3<7>.X 0 0.0749491f
c_82161 XI2.XI1.XI13.XI3<6>.Y 0 0.101266f
c_82179 XI2.XI1.XI13.XI3<7>.NEN 0 0.0870284f
c_82198 XI2.XI1.XI13.XI3<6>.NEN 0 0.0875326f
c_82211 XI2.XI1.XI13.XI3<5>.X 0 0.0749362f
c_82225 XI2.XI1.XI13.XI3<4>.Y 0 0.100334f
c_82243 XI2.XI1.XI13.XI3<5>.NEN 0 0.0868938f
c_82261 XI2.XI1.XI13.XI3<4>.NEN 0 0.0875193f
c_82277 XI2.XI1.XI13.XI3<10>.X 0 0.0748233f
c_82294 XI2.XI1.XI13.XI3<11>.Y 0 0.101302f
c_82309 XI2.XI1.XI13.XI3<11>.X 0 0.0748016f
c_82325 XI2.XI1.XI13.XI3<10>.Y 0 0.101242f
c_82344 XI2.XI1.XI13.XI3<11>.NEN 0 0.0871723f
c_82362 XI2.XI1.XI13.XI3<10>.NEN 0 0.0875864f
c_82376 XI2.XI1.XI13.XI3<9>.X 0 0.0754531f
c_82392 XI2.XI1.XI13.XI3<8>.Y 0 0.101071f
c_82411 XI2.XI1.XI13.XI3<9>.NEN 0 0.0869866f
c_82430 XI2.XI1.XI13.XI3<8>.NEN 0 0.0875468f
c_82448 XI2.XI1.XI13.XI3<14>.X 0 0.0723887f
c_82466 XI2.XI1.XI13.XI3<15>.Y 0 0.0999005f
c_82483 XI2.XI1.XI13.XI3<15>.X 0 0.0735237f
c_82502 XI2.XI1.XI13.XI3<14>.Y 0 0.100702f
c_82519 XI2.XI1.XI13.XI3<15>.NEN 0 0.0877089f
c_82539 XI2.XI1.XI13.XI3<14>.NEN 0 0.0875754f
c_82555 XI2.XI1.XI13.XI3<13>.X 0 0.0737014f
c_82573 XI2.XI1.XI13.XI3<12>.Y 0 0.101125f
c_82593 XI2.XI1.XI13.XI3<13>.NEN 0 0.0869316f
c_82612 XI2.XI1.XI13.XI3<12>.NEN 0 0.0877414f
c_82650 XI1.XI1.WR_EN_BAR 0 2.6598f
c_82657 XI1.XI1.DEC_ADDR_BAR<12> 0 0.130936f
c_82664 XI1.XI1.DEC_ADDR_BAR<11> 0 0.132399f
c_82672 XI1.XI1.DEC_ADDR_BAR<10> 0 0.132579f
c_82680 XI1.XI1.DEC_ADDR_BAR<9> 0 0.132712f
c_82689 XI1.XI1.DEC_ADDR_BAR<8> 0 0.133506f
c_82697 XI1.XI1.DEC_ADDR_BAR<7> 0 0.13353f
c_82707 XI1.XI1.DEC_ADDR_BAR<6> 0 0.132864f
c_82715 XI1.XI1.DEC_ADDR_BAR<5> 0 0.134987f
c_82724 XI1.XI1.DEC_ADDR_BAR<4> 0 0.133506f
c_82732 XI1.XI1.DEC_ADDR_BAR<3> 0 0.13353f
c_82740 XI1.XI1.DEC_ADDR_BAR<2> 0 0.133189f
c_82747 XI1.XI1.DEC_ADDR_BAR<1> 0 0.133568f
c_82754 XI1.XI1.DEC_ADDR_BAR<0> 0 0.136974f
c_82876 XI1.WR_ADDR_EN<12> 0 0.464123f
c_82998 XI1.WR_ADDR_EN<11> 0 0.466512f
c_83120 XI1.WR_ADDR_EN<10> 0 0.465607f
c_83242 XI1.WR_ADDR_EN<9> 0 0.466512f
c_83364 XI1.WR_ADDR_EN<8> 0 0.466512f
c_83486 XI1.WR_ADDR_EN<7> 0 0.466512f
c_83608 XI1.WR_ADDR_EN<6> 0 0.460705f
c_83730 XI1.WR_ADDR_EN<5> 0 0.579683f
c_83852 XI1.WR_ADDR_EN<4> 0 0.58035f
c_83974 XI1.WR_ADDR_EN<3> 0 0.580631f
c_84096 XI1.WR_ADDR_EN<2> 0 0.576248f
c_84218 XI1.WR_ADDR_EN<1> 0 0.576248f
c_84322 XI1.WR_ADDR_EN<0> 0 0.578701f
c_84537 XI1.XI0.CK_EN<12> 0 2.03469f
c_84546 XI1.XI1.XI0.NET_11XX 0 0.15351f
c_84578 XI1.XI1.XI0.NET_XX00 0 1.10672f
c_84602 XI1.XI1.XI0.NET_XX11 0 0.706648f
c_84620 XI1.XI1.XI0.NET_10XX 0 0.635549f
c_84637 XI1.XI1.XI0.ADDR_BAR<2> 0 0.648385f
c_84655 XI1.XI1.XI0.ADDR_BAR<0> 0 0.707917f
c_84681 XI1.XI1.XI0.NET_XX10 0 0.980681f
c_84700 XI1.XI1.XI0.NET_01XX 0 0.611358f
c_84715 XI1.XI1.XI0.ADDR_BAR<1> 0 0.524568f
c_84738 XI1.XI1.XI0.NET_XX01 0 0.970973f
c_84756 XI1.XI1.XI0.NET_00XX 0 0.628192f
c_84773 XI1.XI1.XI0.ADDR_BAR<3> 0 0.394208f
c_84780 XI1.XI1.XI0.XI11.ZN_NEG 0 0.105781f
c_84788 XI1.XI1.XI0.XI7.ZN_NEG 0 0.106313f
c_84797 XI1.XI1.XI0.XI10.ZN_NEG 0 0.105708f
c_84806 XI1.XI1.XI0.XI6.ZN_NEG 0 0.105776f
c_84816 XI1.XI1.XI0.XI9.ZN_NEG 0 0.105064f
c_84826 XI1.XI1.XI0.XI5.ZN_NEG 0 0.105802f
c_84834 XI1.XI1.XI0.XI8.ZN_NEG 0 0.108226f
c_84841 XI1.XI1.XI0.XI4.ZN_NEG 0 0.106004f
c_84977 XI1.XI0.M_DATA<0> 0 1.27533f
c_85099 XI1.XI0.M_DATA<1> 0 1.25318f
c_85222 XI1.XI0.M_DATA<2> 0 1.30822f
c_85335 XI1.XI0.M_DATA<3> 0 1.24773f
c_85446 XI1.XI0.M_DATA<4> 0 1.31264f
c_85547 XI1.XI0.M_DATA<5> 0 1.25623f
c_85645 XI1.XI0.M_DATA<6> 0 1.32522f
c_85743 XI1.XI0.M_DATA<7> 0 1.28923f
c_85854 XI1.XI0.M_DATA<8> 0 1.3155f
c_85964 XI1.XI0.M_DATA<9> 0 1.23728f
c_86063 XI1.XI0.M_DATA<10> 0 1.3873f
c_86161 XI1.XI0.M_DATA<11> 0 1.23697f
c_86272 XI1.XI0.M_DATA<12> 0 1.42212f
c_86382 XI1.XI0.M_DATA<13> 0 1.25778f
c_86506 XI1.XI0.M_DATA<14> 0 1.30028f
c_86628 XI1.XI0.M_DATA<15> 0 1.26199f
c_86768 XI1.XI0.CK 0 2.74687f
c_86996 XI1.XI0.CK_EN<11> 0 1.62067f
c_87225 XI1.XI0.CK_EN<10> 0 1.64196f
c_87453 XI1.XI0.CK_EN<9> 0 1.60463f
c_87682 XI1.XI0.CK_EN<8> 0 1.58805f
c_87911 XI1.XI0.CK_EN<7> 0 1.57509f
c_88142 XI1.XI0.CK_EN<6> 0 1.46249f
c_88368 XI1.XI0.CK_EN<3> 0 1.62261f
c_88398 XI1.XI0.NET18 0 0.182687f
c_88624 XI1.XI0.CLK_N 0 3.22412f
c_88850 XI1.XI0.CK_EN<2> 0 1.89678f
c_88864 XI1.XI0.CLK_PREBUFF 0 0.125876f
c_88882 XI1.XI0.NET5 0 0.0965063f
c_89106 XI1.XI0.CK_EN<1> 0 1.59852f
c_89330 XI1.XI0.CK_EN<0> 0 1.61714f
c_89349 XI1.XI0.NET9 0 0.141401f
c_89364 XI1.XI0.NET13 0 0.0923249f
c_89586 XI1.XI0.CK_EN<5> 0 1.85243f
c_89809 XI1.XI0.CK_EN<4> 0 1.87374f
c_89819 XI1.XI0.XI14<12>.NET_002 0 0.0891143f
c_89827 XI1.XI0.XI14<12>.NET_004 0 0.102508f
c_89838 XI1.XI0.XI14<12>.NET_005 0 0.16956f
c_89855 XI1.XI0.XI14<12>.NET_000 0 0.154126f
c_89867 XI1.XI0.XI14<12>.NET_006 0 0.151967f
c_89877 XI1.XI0.XI14<11>.NET_002 0 0.0853665f
c_89885 XI1.XI0.XI14<11>.NET_004 0 0.100509f
c_89896 XI1.XI0.XI14<11>.NET_005 0 0.169521f
c_89914 XI1.XI0.XI14<11>.NET_000 0 0.153851f
c_89927 XI1.XI0.XI14<11>.NET_006 0 0.14249f
c_89937 XI1.XI0.XI14<10>.NET_002 0 0.0853665f
c_89945 XI1.XI0.XI14<10>.NET_004 0 0.100509f
c_89956 XI1.XI0.XI14<10>.NET_005 0 0.169521f
c_89974 XI1.XI0.XI14<10>.NET_000 0 0.153851f
c_89987 XI1.XI0.XI14<10>.NET_006 0 0.142495f
c_89997 XI1.XI0.XI14<9>.NET_002 0 0.0853665f
c_90005 XI1.XI0.XI14<9>.NET_004 0 0.100509f
c_90016 XI1.XI0.XI14<9>.NET_005 0 0.169521f
c_90034 XI1.XI0.XI14<9>.NET_000 0 0.153827f
c_90047 XI1.XI0.XI14<9>.NET_006 0 0.142495f
c_90057 XI1.XI0.XI14<8>.NET_002 0 0.0853665f
c_90065 XI1.XI0.XI14<8>.NET_004 0 0.100509f
c_90076 XI1.XI0.XI14<8>.NET_005 0 0.169521f
c_90094 XI1.XI0.XI14<8>.NET_000 0 0.153817f
c_90107 XI1.XI0.XI14<8>.NET_006 0 0.142495f
c_90117 XI1.XI0.XI14<7>.NET_002 0 0.0853665f
c_90125 XI1.XI0.XI14<7>.NET_004 0 0.100509f
c_90136 XI1.XI0.XI14<7>.NET_005 0 0.169521f
c_90154 XI1.XI0.XI14<7>.NET_000 0 0.153777f
c_90167 XI1.XI0.XI14<7>.NET_006 0 0.142495f
c_90177 XI1.XI0.XI14<6>.NET_002 0 0.0848409f
c_90185 XI1.XI0.XI14<6>.NET_004 0 0.0972279f
c_90196 XI1.XI0.XI14<6>.NET_005 0 0.168947f
c_90214 XI1.XI0.XI14<6>.NET_000 0 0.152643f
c_90227 XI1.XI0.XI14<6>.NET_006 0 0.142483f
c_90237 XI1.XI0.XI14<5>.NET_002 0 0.0855551f
c_90245 XI1.XI0.XI14<5>.NET_004 0 0.100254f
c_90255 XI1.XI0.XI14<5>.NET_005 0 0.168988f
c_90271 XI1.XI0.XI14<5>.NET_000 0 0.151925f
c_90283 XI1.XI0.XI14<5>.NET_006 0 0.141815f
c_90293 XI1.XI0.XI14<4>.NET_002 0 0.0855551f
c_90301 XI1.XI0.XI14<4>.NET_004 0 0.100509f
c_90311 XI1.XI0.XI14<4>.NET_005 0 0.169495f
c_90327 XI1.XI0.XI14<4>.NET_000 0 0.153851f
c_90339 XI1.XI0.XI14<4>.NET_006 0 0.142312f
c_90349 XI1.XI0.XI14<3>.NET_002 0 0.0855551f
c_90357 XI1.XI0.XI14<3>.NET_004 0 0.100509f
c_90368 XI1.XI0.XI14<3>.NET_005 0 0.169495f
c_90385 XI1.XI0.XI14<3>.NET_000 0 0.153851f
c_90398 XI1.XI0.XI14<3>.NET_006 0 0.142312f
c_90408 XI1.XI0.XI14<2>.NET_002 0 0.0855551f
c_90416 XI1.XI0.XI14<2>.NET_004 0 0.100509f
c_90427 XI1.XI0.XI14<2>.NET_005 0 0.169495f
c_90444 XI1.XI0.XI14<2>.NET_000 0 0.153851f
c_90457 XI1.XI0.XI14<2>.NET_006 0 0.142312f
c_90467 XI1.XI0.XI14<1>.NET_002 0 0.0855551f
c_90475 XI1.XI0.XI14<1>.NET_004 0 0.100509f
c_90486 XI1.XI0.XI14<1>.NET_005 0 0.169495f
c_90503 XI1.XI0.XI14<1>.NET_000 0 0.153851f
c_90516 XI1.XI0.XI14<1>.NET_006 0 0.142312f
c_90525 XI1.XI0.XI14<0>.NET_002 0 0.0851332f
c_90534 XI1.XI0.XI14<0>.NET_004 0 0.100817f
c_90545 XI1.XI0.XI14<0>.NET_005 0 0.170101f
c_90565 XI1.XI0.XI14<0>.NET_000 0 0.171267f
c_90578 XI1.XI0.XI14<0>.NET_006 0 0.142312f
c_90602 XI1.XI0.XI1<12>.XI7<3>.NET_000 0 0.191538f
c_90619 XI1.XI0.XI1<12>.XI7<3>.NET_001 0 0.068031f
c_90637 XI1.XI0.XI1<12>.XI7<3>.NET_003 0 0.182225f
c_90652 XI1.XI0.XI1<12>.XI7<3>.NET_005 0 0.0724441f
c_90673 XI1.XI0.XI1<12>.XI7<2>.NET_000 0 0.190975f
c_90691 XI1.XI0.XI1<12>.XI7<2>.NET_001 0 0.0660846f
c_90711 XI1.XI0.XI1<12>.XI7<2>.NET_003 0 0.181683f
c_90726 XI1.XI0.XI1<12>.XI7<2>.NET_005 0 0.0724441f
c_90748 XI1.XI0.XI1<12>.XI7<1>.NET_000 0 0.190139f
c_90765 XI1.XI0.XI1<12>.XI7<1>.NET_001 0 0.0675987f
c_90783 XI1.XI0.XI1<12>.XI7<1>.NET_003 0 0.182438f
c_90798 XI1.XI0.XI1<12>.XI7<1>.NET_005 0 0.0724441f
c_90819 XI1.XI0.XI1<12>.XI7<0>.NET_000 0 0.192932f
c_90835 XI1.XI0.XI1<12>.XI7<0>.NET_001 0 0.0661732f
c_90854 XI1.XI0.XI1<12>.XI7<0>.NET_003 0 0.183265f
c_90870 XI1.XI0.XI1<12>.XI7<0>.NET_005 0 0.0724585f
c_90887 XI1.XI0.XI1<12>.XI7<7>.NET_000 0 0.200287f
c_90903 XI1.XI0.XI1<12>.XI7<7>.NET_001 0 0.0680598f
c_90919 XI1.XI0.XI1<12>.XI7<7>.NET_003 0 0.184508f
c_90934 XI1.XI0.XI1<12>.XI7<7>.NET_005 0 0.0723879f
c_90956 XI1.XI0.XI1<12>.XI7<6>.NET_000 0 0.194467f
c_90973 XI1.XI0.XI1<12>.XI7<6>.NET_001 0 0.0662675f
c_90991 XI1.XI0.XI1<12>.XI7<6>.NET_003 0 0.182351f
c_91006 XI1.XI0.XI1<12>.XI7<6>.NET_005 0 0.0724441f
c_91031 XI1.XI0.XI1<12>.XI7<5>.NET_000 0 0.186674f
c_91047 XI1.XI0.XI1<12>.XI7<5>.NET_001 0 0.0673432f
c_91065 XI1.XI0.XI1<12>.XI7<5>.NET_003 0 0.182836f
c_91080 XI1.XI0.XI1<12>.XI7<5>.NET_005 0 0.0724441f
c_91105 XI1.XI0.XI1<12>.XI7<4>.NET_000 0 0.187092f
c_91122 XI1.XI0.XI1<12>.XI7<4>.NET_001 0 0.0667151f
c_91141 XI1.XI0.XI1<12>.XI7<4>.NET_003 0 0.18174f
c_91156 XI1.XI0.XI1<12>.XI7<4>.NET_005 0 0.0724441f
c_91176 XI1.XI0.XI1<12>.XI7<11>.NET_000 0 0.19187f
c_91192 XI1.XI0.XI1<12>.XI7<11>.NET_001 0 0.0681178f
c_91209 XI1.XI0.XI1<12>.XI7<11>.NET_003 0 0.183007f
c_91225 XI1.XI0.XI1<12>.XI7<11>.NET_005 0 0.0724441f
c_91245 XI1.XI0.XI1<12>.XI7<10>.NET_000 0 0.19353f
c_91260 XI1.XI0.XI1<12>.XI7<10>.NET_001 0 0.0662224f
c_91276 XI1.XI0.XI1<12>.XI7<10>.NET_003 0 0.183599f
c_91292 XI1.XI0.XI1<12>.XI7<10>.NET_005 0 0.0724441f
c_91311 XI1.XI0.XI1<12>.XI7<9>.NET_000 0 0.192221f
c_91328 XI1.XI0.XI1<12>.XI7<9>.NET_001 0 0.0678273f
c_91346 XI1.XI0.XI1<12>.XI7<9>.NET_003 0 0.182748f
c_91362 XI1.XI0.XI1<12>.XI7<9>.NET_005 0 0.0724441f
c_91383 XI1.XI0.XI1<12>.XI7<8>.NET_000 0 0.198921f
c_91400 XI1.XI0.XI1<12>.XI7<8>.NET_001 0 0.0659516f
c_91418 XI1.XI0.XI1<12>.XI7<8>.NET_003 0 0.182267f
c_91434 XI1.XI0.XI1<12>.XI7<8>.NET_005 0 0.0721711f
c_91455 XI1.XI0.XI1<12>.XI7<15>.NET_000 0 0.186734f
c_91473 XI1.XI0.XI1<12>.XI7<15>.NET_001 0 0.0681481f
c_91491 XI1.XI0.XI1<12>.XI7<15>.NET_003 0 0.183371f
c_91507 XI1.XI0.XI1<12>.XI7<15>.NET_005 0 0.0727082f
c_91527 XI1.XI0.XI1<12>.XI7<14>.NET_000 0 0.190158f
c_91544 XI1.XI0.XI1<12>.XI7<14>.NET_001 0 0.0658913f
c_91562 XI1.XI0.XI1<12>.XI7<14>.NET_003 0 0.182032f
c_91578 XI1.XI0.XI1<12>.XI7<14>.NET_005 0 0.0724441f
c_91600 XI1.XI0.XI1<12>.XI7<13>.NET_000 0 0.190435f
c_91617 XI1.XI0.XI1<12>.XI7<13>.NET_001 0 0.0687736f
c_91635 XI1.XI0.XI1<12>.XI7<13>.NET_003 0 0.183668f
c_91651 XI1.XI0.XI1<12>.XI7<13>.NET_005 0 0.0724835f
c_91671 XI1.XI0.XI1<12>.XI7<12>.NET_000 0 0.19446f
c_91686 XI1.XI0.XI1<12>.XI7<12>.NET_001 0 0.0658629f
c_91702 XI1.XI0.XI1<12>.XI7<12>.NET_003 0 0.185262f
c_91717 XI1.XI0.XI1<12>.XI7<12>.NET_005 0 0.0732094f
c_91738 XI1.XI0.XI1<11>.XI7<3>.NET_000 0 0.187398f
c_91755 XI1.XI0.XI1<11>.XI7<3>.NET_001 0 0.0680399f
c_91773 XI1.XI0.XI1<11>.XI7<3>.NET_003 0 0.181695f
c_91788 XI1.XI0.XI1<11>.XI7<3>.NET_005 0 0.0724441f
c_91810 XI1.XI0.XI1<11>.XI7<2>.NET_000 0 0.187414f
c_91828 XI1.XI0.XI1<11>.XI7<2>.NET_001 0 0.0671465f
c_91848 XI1.XI0.XI1<11>.XI7<2>.NET_003 0 0.180896f
c_91863 XI1.XI0.XI1<11>.XI7<2>.NET_005 0 0.0724441f
c_91884 XI1.XI0.XI1<11>.XI7<1>.NET_000 0 0.186653f
c_91901 XI1.XI0.XI1<11>.XI7<1>.NET_001 0 0.0676071f
c_91919 XI1.XI0.XI1<11>.XI7<1>.NET_003 0 0.181903f
c_91934 XI1.XI0.XI1<11>.XI7<1>.NET_005 0 0.0724441f
c_91956 XI1.XI0.XI1<11>.XI7<0>.NET_000 0 0.191214f
c_91973 XI1.XI0.XI1<11>.XI7<0>.NET_001 0 0.0671299f
c_91992 XI1.XI0.XI1<11>.XI7<0>.NET_003 0 0.182475f
c_92008 XI1.XI0.XI1<11>.XI7<0>.NET_005 0 0.0724585f
c_92026 XI1.XI0.XI1<11>.XI7<7>.NET_000 0 0.197474f
c_92042 XI1.XI0.XI1<11>.XI7<7>.NET_001 0 0.0677901f
c_92058 XI1.XI0.XI1<11>.XI7<7>.NET_003 0 0.183947f
c_92073 XI1.XI0.XI1<11>.XI7<7>.NET_005 0 0.0723879f
c_92093 XI1.XI0.XI1<11>.XI7<6>.NET_000 0 0.189436f
c_92110 XI1.XI0.XI1<11>.XI7<6>.NET_001 0 0.0671634f
c_92128 XI1.XI0.XI1<11>.XI7<6>.NET_003 0 0.181534f
c_92143 XI1.XI0.XI1<11>.XI7<6>.NET_005 0 0.0724441f
c_92163 XI1.XI0.XI1<11>.XI7<5>.NET_000 0 0.18932f
c_92179 XI1.XI0.XI1<11>.XI7<5>.NET_001 0 0.0678117f
c_92197 XI1.XI0.XI1<11>.XI7<5>.NET_003 0 0.182305f
c_92212 XI1.XI0.XI1<11>.XI7<5>.NET_005 0 0.0724441f
c_92233 XI1.XI0.XI1<11>.XI7<4>.NET_000 0 0.18791f
c_92250 XI1.XI0.XI1<11>.XI7<4>.NET_001 0 0.0676945f
c_92269 XI1.XI0.XI1<11>.XI7<4>.NET_003 0 0.180948f
c_92284 XI1.XI0.XI1<11>.XI7<4>.NET_005 0 0.0724441f
c_92304 XI1.XI0.XI1<11>.XI7<11>.NET_000 0 0.189304f
c_92320 XI1.XI0.XI1<11>.XI7<11>.NET_001 0 0.0685193f
c_92337 XI1.XI0.XI1<11>.XI7<11>.NET_003 0 0.182476f
c_92353 XI1.XI0.XI1<11>.XI7<11>.NET_005 0 0.0724441f
c_92372 XI1.XI0.XI1<11>.XI7<10>.NET_000 0 0.190142f
c_92387 XI1.XI0.XI1<11>.XI7<10>.NET_001 0 0.0671183f
c_92403 XI1.XI0.XI1<11>.XI7<10>.NET_003 0 0.182799f
c_92419 XI1.XI0.XI1<11>.XI7<10>.NET_005 0 0.0724441f
c_92440 XI1.XI0.XI1<11>.XI7<9>.NET_000 0 0.18983f
c_92457 XI1.XI0.XI1<11>.XI7<9>.NET_001 0 0.0683151f
c_92475 XI1.XI0.XI1<11>.XI7<9>.NET_003 0 0.18232f
c_92491 XI1.XI0.XI1<11>.XI7<9>.NET_005 0 0.0724441f
c_92513 XI1.XI0.XI1<11>.XI7<8>.NET_000 0 0.195684f
c_92529 XI1.XI0.XI1<11>.XI7<8>.NET_001 0 0.0669071f
c_92546 XI1.XI0.XI1<11>.XI7<8>.NET_003 0 0.181619f
c_92562 XI1.XI0.XI1<11>.XI7<8>.NET_005 0 0.0721711f
c_92583 XI1.XI0.XI1<11>.XI7<15>.NET_000 0 0.190081f
c_92601 XI1.XI0.XI1<11>.XI7<15>.NET_001 0 0.0676928f
c_92619 XI1.XI0.XI1<11>.XI7<15>.NET_003 0 0.182845f
c_92635 XI1.XI0.XI1<11>.XI7<15>.NET_005 0 0.0727082f
c_92656 XI1.XI0.XI1<11>.XI7<14>.NET_000 0 0.187306f
c_92673 XI1.XI0.XI1<11>.XI7<14>.NET_001 0 0.0669713f
c_92691 XI1.XI0.XI1<11>.XI7<14>.NET_003 0 0.181234f
c_92707 XI1.XI0.XI1<11>.XI7<14>.NET_005 0 0.0724441f
c_92728 XI1.XI0.XI1<11>.XI7<13>.NET_000 0 0.18825f
c_92745 XI1.XI0.XI1<11>.XI7<13>.NET_001 0 0.0689289f
c_92763 XI1.XI0.XI1<11>.XI7<13>.NET_003 0 0.183155f
c_92779 XI1.XI0.XI1<11>.XI7<13>.NET_005 0 0.0724835f
c_92798 XI1.XI0.XI1<11>.XI7<12>.NET_000 0 0.191272f
c_92813 XI1.XI0.XI1<11>.XI7<12>.NET_001 0 0.0667363f
c_92829 XI1.XI0.XI1<11>.XI7<12>.NET_003 0 0.184465f
c_92844 XI1.XI0.XI1<11>.XI7<12>.NET_005 0 0.0732094f
c_92865 XI1.XI0.XI1<10>.XI7<3>.NET_000 0 0.187398f
c_92882 XI1.XI0.XI1<10>.XI7<3>.NET_001 0 0.0680399f
c_92900 XI1.XI0.XI1<10>.XI7<3>.NET_003 0 0.181695f
c_92915 XI1.XI0.XI1<10>.XI7<3>.NET_005 0 0.0724441f
c_92937 XI1.XI0.XI1<10>.XI7<2>.NET_000 0 0.187429f
c_92955 XI1.XI0.XI1<10>.XI7<2>.NET_001 0 0.0671614f
c_92975 XI1.XI0.XI1<10>.XI7<2>.NET_003 0 0.180902f
c_92990 XI1.XI0.XI1<10>.XI7<2>.NET_005 0 0.0724441f
c_93011 XI1.XI0.XI1<10>.XI7<1>.NET_000 0 0.186653f
c_93028 XI1.XI0.XI1<10>.XI7<1>.NET_001 0 0.0676071f
c_93046 XI1.XI0.XI1<10>.XI7<1>.NET_003 0 0.181903f
c_93061 XI1.XI0.XI1<10>.XI7<1>.NET_005 0 0.0724441f
c_93083 XI1.XI0.XI1<10>.XI7<0>.NET_000 0 0.191315f
c_93100 XI1.XI0.XI1<10>.XI7<0>.NET_001 0 0.0671766f
c_93119 XI1.XI0.XI1<10>.XI7<0>.NET_003 0 0.182479f
c_93135 XI1.XI0.XI1<10>.XI7<0>.NET_005 0 0.0724585f
c_93153 XI1.XI0.XI1<10>.XI7<7>.NET_000 0 0.197474f
c_93169 XI1.XI0.XI1<10>.XI7<7>.NET_001 0 0.0677901f
c_93185 XI1.XI0.XI1<10>.XI7<7>.NET_003 0 0.183947f
c_93200 XI1.XI0.XI1<10>.XI7<7>.NET_005 0 0.072441f
c_93220 XI1.XI0.XI1<10>.XI7<6>.NET_000 0 0.18943f
c_93237 XI1.XI0.XI1<10>.XI7<6>.NET_001 0 0.0671634f
c_93255 XI1.XI0.XI1<10>.XI7<6>.NET_003 0 0.181513f
c_93270 XI1.XI0.XI1<10>.XI7<6>.NET_005 0 0.0724441f
c_93290 XI1.XI0.XI1<10>.XI7<5>.NET_000 0 0.18932f
c_93306 XI1.XI0.XI1<10>.XI7<5>.NET_001 0 0.0678117f
c_93324 XI1.XI0.XI1<10>.XI7<5>.NET_003 0 0.182305f
c_93339 XI1.XI0.XI1<10>.XI7<5>.NET_005 0 0.0724441f
c_93360 XI1.XI0.XI1<10>.XI7<4>.NET_000 0 0.18791f
c_93377 XI1.XI0.XI1<10>.XI7<4>.NET_001 0 0.0676945f
c_93396 XI1.XI0.XI1<10>.XI7<4>.NET_003 0 0.180928f
c_93411 XI1.XI0.XI1<10>.XI7<4>.NET_005 0 0.0724441f
c_93431 XI1.XI0.XI1<10>.XI7<11>.NET_000 0 0.189304f
c_93447 XI1.XI0.XI1<10>.XI7<11>.NET_001 0 0.0685193f
c_93464 XI1.XI0.XI1<10>.XI7<11>.NET_003 0 0.182476f
c_93480 XI1.XI0.XI1<10>.XI7<11>.NET_005 0 0.0724441f
c_93499 XI1.XI0.XI1<10>.XI7<10>.NET_000 0 0.190142f
c_93514 XI1.XI0.XI1<10>.XI7<10>.NET_001 0 0.0671183f
c_93530 XI1.XI0.XI1<10>.XI7<10>.NET_003 0 0.182799f
c_93546 XI1.XI0.XI1<10>.XI7<10>.NET_005 0 0.0724441f
c_93567 XI1.XI0.XI1<10>.XI7<9>.NET_000 0 0.189836f
c_93584 XI1.XI0.XI1<10>.XI7<9>.NET_001 0 0.0683151f
c_93602 XI1.XI0.XI1<10>.XI7<9>.NET_003 0 0.182342f
c_93618 XI1.XI0.XI1<10>.XI7<9>.NET_005 0 0.0724441f
c_93640 XI1.XI0.XI1<10>.XI7<8>.NET_000 0 0.195684f
c_93656 XI1.XI0.XI1<10>.XI7<8>.NET_001 0 0.0669071f
c_93673 XI1.XI0.XI1<10>.XI7<8>.NET_003 0 0.181619f
c_93689 XI1.XI0.XI1<10>.XI7<8>.NET_005 0 0.0721711f
c_93710 XI1.XI0.XI1<10>.XI7<15>.NET_000 0 0.190042f
c_93728 XI1.XI0.XI1<10>.XI7<15>.NET_001 0 0.0676565f
c_93746 XI1.XI0.XI1<10>.XI7<15>.NET_003 0 0.182845f
c_93762 XI1.XI0.XI1<10>.XI7<15>.NET_005 0 0.0727082f
c_93783 XI1.XI0.XI1<10>.XI7<14>.NET_000 0 0.187306f
c_93800 XI1.XI0.XI1<10>.XI7<14>.NET_001 0 0.0669713f
c_93818 XI1.XI0.XI1<10>.XI7<14>.NET_003 0 0.181234f
c_93834 XI1.XI0.XI1<10>.XI7<14>.NET_005 0 0.0724441f
c_93855 XI1.XI0.XI1<10>.XI7<13>.NET_000 0 0.18825f
c_93872 XI1.XI0.XI1<10>.XI7<13>.NET_001 0 0.0689289f
c_93890 XI1.XI0.XI1<10>.XI7<13>.NET_003 0 0.183155f
c_93906 XI1.XI0.XI1<10>.XI7<13>.NET_005 0 0.0724835f
c_93925 XI1.XI0.XI1<10>.XI7<12>.NET_000 0 0.191272f
c_93940 XI1.XI0.XI1<10>.XI7<12>.NET_001 0 0.0667363f
c_93956 XI1.XI0.XI1<10>.XI7<12>.NET_003 0 0.184465f
c_93971 XI1.XI0.XI1<10>.XI7<12>.NET_005 0 0.0732094f
c_93992 XI1.XI0.XI1<9>.XI7<3>.NET_000 0 0.187398f
c_94009 XI1.XI0.XI1<9>.XI7<3>.NET_001 0 0.0680399f
c_94027 XI1.XI0.XI1<9>.XI7<3>.NET_003 0 0.181695f
c_94042 XI1.XI0.XI1<9>.XI7<3>.NET_005 0 0.0724441f
c_94064 XI1.XI0.XI1<9>.XI7<2>.NET_000 0 0.187429f
c_94082 XI1.XI0.XI1<9>.XI7<2>.NET_001 0 0.0671614f
c_94102 XI1.XI0.XI1<9>.XI7<2>.NET_003 0 0.180882f
c_94117 XI1.XI0.XI1<9>.XI7<2>.NET_005 0 0.0724441f
c_94138 XI1.XI0.XI1<9>.XI7<1>.NET_000 0 0.186653f
c_94155 XI1.XI0.XI1<9>.XI7<1>.NET_001 0 0.0676071f
c_94173 XI1.XI0.XI1<9>.XI7<1>.NET_003 0 0.181903f
c_94188 XI1.XI0.XI1<9>.XI7<1>.NET_005 0 0.0724441f
c_94210 XI1.XI0.XI1<9>.XI7<0>.NET_000 0 0.191351f
c_94227 XI1.XI0.XI1<9>.XI7<0>.NET_001 0 0.0672151f
c_94246 XI1.XI0.XI1<9>.XI7<0>.NET_003 0 0.182485f
c_94262 XI1.XI0.XI1<9>.XI7<0>.NET_005 0 0.0724585f
c_94281 XI1.XI0.XI1<9>.XI7<7>.NET_000 0 0.197706f
c_94298 XI1.XI0.XI1<9>.XI7<7>.NET_001 0 0.0680096f
c_94315 XI1.XI0.XI1<9>.XI7<7>.NET_003 0 0.183824f
c_94330 XI1.XI0.XI1<9>.XI7<7>.NET_005 0 0.072441f
c_94350 XI1.XI0.XI1<9>.XI7<6>.NET_000 0 0.189397f
c_94367 XI1.XI0.XI1<9>.XI7<6>.NET_001 0 0.0671341f
c_94385 XI1.XI0.XI1<9>.XI7<6>.NET_003 0 0.181409f
c_94400 XI1.XI0.XI1<9>.XI7<6>.NET_005 0 0.0724441f
c_94420 XI1.XI0.XI1<9>.XI7<5>.NET_000 0 0.18932f
c_94436 XI1.XI0.XI1<9>.XI7<5>.NET_001 0 0.0678117f
c_94454 XI1.XI0.XI1<9>.XI7<5>.NET_003 0 0.182305f
c_94469 XI1.XI0.XI1<9>.XI7<5>.NET_005 0 0.0724441f
c_94490 XI1.XI0.XI1<9>.XI7<4>.NET_000 0 0.187904f
c_94507 XI1.XI0.XI1<9>.XI7<4>.NET_001 0 0.0676945f
c_94526 XI1.XI0.XI1<9>.XI7<4>.NET_003 0 0.180907f
c_94541 XI1.XI0.XI1<9>.XI7<4>.NET_005 0 0.0724441f
c_94561 XI1.XI0.XI1<9>.XI7<11>.NET_000 0 0.189288f
c_94577 XI1.XI0.XI1<9>.XI7<11>.NET_001 0 0.0685045f
c_94594 XI1.XI0.XI1<9>.XI7<11>.NET_003 0 0.182465f
c_94610 XI1.XI0.XI1<9>.XI7<11>.NET_005 0 0.0724441f
c_94629 XI1.XI0.XI1<9>.XI7<10>.NET_000 0 0.190142f
c_94644 XI1.XI0.XI1<9>.XI7<10>.NET_001 0 0.0671183f
c_94660 XI1.XI0.XI1<9>.XI7<10>.NET_003 0 0.182799f
c_94676 XI1.XI0.XI1<9>.XI7<10>.NET_005 0 0.0724441f
c_94697 XI1.XI0.XI1<9>.XI7<9>.NET_000 0 0.189836f
c_94714 XI1.XI0.XI1<9>.XI7<9>.NET_001 0 0.0683151f
c_94732 XI1.XI0.XI1<9>.XI7<9>.NET_003 0 0.182367f
c_94748 XI1.XI0.XI1<9>.XI7<9>.NET_005 0 0.0724441f
c_94770 XI1.XI0.XI1<9>.XI7<8>.NET_000 0 0.195684f
c_94786 XI1.XI0.XI1<9>.XI7<8>.NET_001 0 0.0669071f
c_94803 XI1.XI0.XI1<9>.XI7<8>.NET_003 0 0.181619f
c_94819 XI1.XI0.XI1<9>.XI7<8>.NET_005 0 0.0721711f
c_94840 XI1.XI0.XI1<9>.XI7<15>.NET_000 0 0.189948f
c_94858 XI1.XI0.XI1<9>.XI7<15>.NET_001 0 0.067619f
c_94876 XI1.XI0.XI1<9>.XI7<15>.NET_003 0 0.182827f
c_94892 XI1.XI0.XI1<9>.XI7<15>.NET_005 0 0.0727082f
c_94913 XI1.XI0.XI1<9>.XI7<14>.NET_000 0 0.187306f
c_94930 XI1.XI0.XI1<9>.XI7<14>.NET_001 0 0.0669713f
c_94948 XI1.XI0.XI1<9>.XI7<14>.NET_003 0 0.181234f
c_94964 XI1.XI0.XI1<9>.XI7<14>.NET_005 0 0.0724441f
c_94985 XI1.XI0.XI1<9>.XI7<13>.NET_000 0 0.188234f
c_95002 XI1.XI0.XI1<9>.XI7<13>.NET_001 0 0.068914f
c_95020 XI1.XI0.XI1<9>.XI7<13>.NET_003 0 0.183144f
c_95036 XI1.XI0.XI1<9>.XI7<13>.NET_005 0 0.0724835f
c_95055 XI1.XI0.XI1<9>.XI7<12>.NET_000 0 0.191272f
c_95070 XI1.XI0.XI1<9>.XI7<12>.NET_001 0 0.0667363f
c_95086 XI1.XI0.XI1<9>.XI7<12>.NET_003 0 0.184465f
c_95101 XI1.XI0.XI1<9>.XI7<12>.NET_005 0 0.0732094f
c_95122 XI1.XI0.XI1<8>.XI7<3>.NET_000 0 0.187398f
c_95139 XI1.XI0.XI1<8>.XI7<3>.NET_001 0 0.0680399f
c_95157 XI1.XI0.XI1<8>.XI7<3>.NET_003 0 0.181695f
c_95172 XI1.XI0.XI1<8>.XI7<3>.NET_005 0 0.0724441f
c_95194 XI1.XI0.XI1<8>.XI7<2>.NET_000 0 0.187421f
c_95212 XI1.XI0.XI1<8>.XI7<2>.NET_001 0 0.0671614f
c_95232 XI1.XI0.XI1<8>.XI7<2>.NET_003 0 0.180861f
c_95247 XI1.XI0.XI1<8>.XI7<2>.NET_005 0 0.0724441f
c_95268 XI1.XI0.XI1<8>.XI7<1>.NET_000 0 0.186653f
c_95285 XI1.XI0.XI1<8>.XI7<1>.NET_001 0 0.0676071f
c_95303 XI1.XI0.XI1<8>.XI7<1>.NET_003 0 0.181903f
c_95318 XI1.XI0.XI1<8>.XI7<1>.NET_005 0 0.0724441f
c_95340 XI1.XI0.XI1<8>.XI7<0>.NET_000 0 0.19136f
c_95357 XI1.XI0.XI1<8>.XI7<0>.NET_001 0 0.0672254f
c_95376 XI1.XI0.XI1<8>.XI7<0>.NET_003 0 0.182465f
c_95392 XI1.XI0.XI1<8>.XI7<0>.NET_005 0 0.0724585f
c_95411 XI1.XI0.XI1<8>.XI7<7>.NET_000 0 0.197752f
c_95428 XI1.XI0.XI1<8>.XI7<7>.NET_001 0 0.0680304f
c_95445 XI1.XI0.XI1<8>.XI7<7>.NET_003 0 0.183961f
c_95460 XI1.XI0.XI1<8>.XI7<7>.NET_005 0 0.0723879f
c_95479 XI1.XI0.XI1<8>.XI7<6>.NET_000 0 0.189436f
c_95495 XI1.XI0.XI1<8>.XI7<6>.NET_001 0 0.0671634f
c_95512 XI1.XI0.XI1<8>.XI7<6>.NET_003 0 0.181559f
c_95527 XI1.XI0.XI1<8>.XI7<6>.NET_005 0 0.0724441f
c_95548 XI1.XI0.XI1<8>.XI7<5>.NET_000 0 0.189281f
c_95565 XI1.XI0.XI1<8>.XI7<5>.NET_001 0 0.0677824f
c_95584 XI1.XI0.XI1<8>.XI7<5>.NET_003 0 0.182156f
c_95599 XI1.XI0.XI1<8>.XI7<5>.NET_005 0 0.0724441f
c_95620 XI1.XI0.XI1<8>.XI7<4>.NET_000 0 0.18787f
c_95637 XI1.XI0.XI1<8>.XI7<4>.NET_001 0 0.0676652f
c_95656 XI1.XI0.XI1<8>.XI7<4>.NET_003 0 0.180803f
c_95671 XI1.XI0.XI1<8>.XI7<4>.NET_005 0 0.0724441f
c_95691 XI1.XI0.XI1<8>.XI7<11>.NET_000 0 0.189268f
c_95707 XI1.XI0.XI1<8>.XI7<11>.NET_001 0 0.0685029f
c_95724 XI1.XI0.XI1<8>.XI7<11>.NET_003 0 0.182455f
c_95740 XI1.XI0.XI1<8>.XI7<11>.NET_005 0 0.0724441f
c_95759 XI1.XI0.XI1<8>.XI7<10>.NET_000 0 0.190142f
c_95774 XI1.XI0.XI1<8>.XI7<10>.NET_001 0 0.0671183f
c_95790 XI1.XI0.XI1<8>.XI7<10>.NET_003 0 0.182799f
c_95806 XI1.XI0.XI1<8>.XI7<10>.NET_005 0 0.0724441f
c_95827 XI1.XI0.XI1<8>.XI7<9>.NET_000 0 0.18982f
c_95844 XI1.XI0.XI1<8>.XI7<9>.NET_001 0 0.0683002f
c_95862 XI1.XI0.XI1<8>.XI7<9>.NET_003 0 0.182356f
c_95878 XI1.XI0.XI1<8>.XI7<9>.NET_005 0 0.0724441f
c_95900 XI1.XI0.XI1<8>.XI7<8>.NET_000 0 0.195684f
c_95916 XI1.XI0.XI1<8>.XI7<8>.NET_001 0 0.0669071f
c_95933 XI1.XI0.XI1<8>.XI7<8>.NET_003 0 0.181619f
c_95949 XI1.XI0.XI1<8>.XI7<8>.NET_005 0 0.0721711f
c_95969 XI1.XI0.XI1<8>.XI7<15>.NET_000 0 0.190105f
c_95986 XI1.XI0.XI1<8>.XI7<15>.NET_001 0 0.0677275f
c_96004 XI1.XI0.XI1<8>.XI7<15>.NET_003 0 0.18282f
c_96020 XI1.XI0.XI1<8>.XI7<15>.NET_005 0 0.0727082f
c_96041 XI1.XI0.XI1<8>.XI7<14>.NET_000 0 0.187306f
c_96058 XI1.XI0.XI1<8>.XI7<14>.NET_001 0 0.0669713f
c_96076 XI1.XI0.XI1<8>.XI7<14>.NET_003 0 0.181234f
c_96092 XI1.XI0.XI1<8>.XI7<14>.NET_005 0 0.0724441f
c_96113 XI1.XI0.XI1<8>.XI7<13>.NET_000 0 0.188213f
c_96130 XI1.XI0.XI1<8>.XI7<13>.NET_001 0 0.0689125f
c_96148 XI1.XI0.XI1<8>.XI7<13>.NET_003 0 0.183134f
c_96164 XI1.XI0.XI1<8>.XI7<13>.NET_005 0 0.0724835f
c_96183 XI1.XI0.XI1<8>.XI7<12>.NET_000 0 0.191272f
c_96198 XI1.XI0.XI1<8>.XI7<12>.NET_001 0 0.0667363f
c_96214 XI1.XI0.XI1<8>.XI7<12>.NET_003 0 0.184465f
c_96229 XI1.XI0.XI1<8>.XI7<12>.NET_005 0 0.0732094f
c_96251 XI1.XI0.XI1<7>.XI7<3>.NET_000 0 0.187359f
c_96269 XI1.XI0.XI1<7>.XI7<3>.NET_001 0 0.0680097f
c_96288 XI1.XI0.XI1<7>.XI7<3>.NET_003 0 0.181545f
c_96303 XI1.XI0.XI1<7>.XI7<3>.NET_005 0 0.0724441f
c_96325 XI1.XI0.XI1<7>.XI7<2>.NET_000 0 0.18739f
c_96343 XI1.XI0.XI1<7>.XI7<2>.NET_001 0 0.0671614f
c_96363 XI1.XI0.XI1<7>.XI7<2>.NET_003 0 0.180758f
c_96378 XI1.XI0.XI1<7>.XI7<2>.NET_005 0 0.0724441f
c_96399 XI1.XI0.XI1<7>.XI7<1>.NET_000 0 0.186653f
c_96416 XI1.XI0.XI1<7>.XI7<1>.NET_001 0 0.0676071f
c_96434 XI1.XI0.XI1<7>.XI7<1>.NET_003 0 0.181903f
c_96449 XI1.XI0.XI1<7>.XI7<1>.NET_005 0 0.0724441f
c_96471 XI1.XI0.XI1<7>.XI7<0>.NET_000 0 0.191358f
c_96488 XI1.XI0.XI1<7>.XI7<0>.NET_001 0 0.0672319f
c_96507 XI1.XI0.XI1<7>.XI7<0>.NET_003 0 0.182443f
c_96523 XI1.XI0.XI1<7>.XI7<0>.NET_005 0 0.0724585f
c_96542 XI1.XI0.XI1<7>.XI7<7>.NET_000 0 0.197691f
c_96559 XI1.XI0.XI1<7>.XI7<7>.NET_001 0 0.0680461f
c_96576 XI1.XI0.XI1<7>.XI7<7>.NET_003 0 0.183947f
c_96591 XI1.XI0.XI1<7>.XI7<7>.NET_005 0 0.0723879f
c_96610 XI1.XI0.XI1<7>.XI7<6>.NET_000 0 0.189436f
c_96626 XI1.XI0.XI1<7>.XI7<6>.NET_001 0 0.0671634f
c_96643 XI1.XI0.XI1<7>.XI7<6>.NET_003 0 0.181559f
c_96658 XI1.XI0.XI1<7>.XI7<6>.NET_005 0 0.0724441f
c_96679 XI1.XI0.XI1<7>.XI7<5>.NET_000 0 0.189314f
c_96696 XI1.XI0.XI1<7>.XI7<5>.NET_001 0 0.0678117f
c_96715 XI1.XI0.XI1<7>.XI7<5>.NET_003 0 0.182259f
c_96730 XI1.XI0.XI1<7>.XI7<5>.NET_005 0 0.0724441f
c_96750 XI1.XI0.XI1<7>.XI7<4>.NET_000 0 0.18791f
c_96766 XI1.XI0.XI1<7>.XI7<4>.NET_001 0 0.0676945f
c_96784 XI1.XI0.XI1<7>.XI7<4>.NET_003 0 0.180953f
c_96799 XI1.XI0.XI1<7>.XI7<4>.NET_005 0 0.0724441f
c_96818 XI1.XI0.XI1<7>.XI7<11>.NET_000 0 0.189304f
c_96833 XI1.XI0.XI1<7>.XI7<11>.NET_001 0 0.0685193f
c_96850 XI1.XI0.XI1<7>.XI7<11>.NET_003 0 0.182449f
c_96866 XI1.XI0.XI1<7>.XI7<11>.NET_005 0 0.0724441f
c_96885 XI1.XI0.XI1<7>.XI7<10>.NET_000 0 0.190142f
c_96900 XI1.XI0.XI1<7>.XI7<10>.NET_001 0 0.0671183f
c_96916 XI1.XI0.XI1<7>.XI7<10>.NET_003 0 0.182799f
c_96932 XI1.XI0.XI1<7>.XI7<10>.NET_005 0 0.0724441f
c_96953 XI1.XI0.XI1<7>.XI7<9>.NET_000 0 0.1898f
c_96970 XI1.XI0.XI1<7>.XI7<9>.NET_001 0 0.0682986f
c_96988 XI1.XI0.XI1<7>.XI7<9>.NET_003 0 0.182345f
c_97004 XI1.XI0.XI1<7>.XI7<9>.NET_005 0 0.0724441f
c_97026 XI1.XI0.XI1<7>.XI7<8>.NET_000 0 0.195684f
c_97042 XI1.XI0.XI1<7>.XI7<8>.NET_001 0 0.0669071f
c_97059 XI1.XI0.XI1<7>.XI7<8>.NET_003 0 0.181619f
c_97075 XI1.XI0.XI1<7>.XI7<8>.NET_005 0 0.0721711f
c_97095 XI1.XI0.XI1<7>.XI7<15>.NET_000 0 0.190105f
c_97112 XI1.XI0.XI1<7>.XI7<15>.NET_001 0 0.0677275f
c_97129 XI1.XI0.XI1<7>.XI7<15>.NET_003 0 0.182845f
c_97145 XI1.XI0.XI1<7>.XI7<15>.NET_005 0 0.0727082f
c_97166 XI1.XI0.XI1<7>.XI7<14>.NET_000 0 0.187306f
c_97183 XI1.XI0.XI1<7>.XI7<14>.NET_001 0 0.0669713f
c_97202 XI1.XI0.XI1<7>.XI7<14>.NET_003 0 0.181207f
c_97218 XI1.XI0.XI1<7>.XI7<14>.NET_005 0 0.0724441f
c_97238 XI1.XI0.XI1<7>.XI7<13>.NET_000 0 0.18825f
c_97254 XI1.XI0.XI1<7>.XI7<13>.NET_001 0 0.0689289f
c_97272 XI1.XI0.XI1<7>.XI7<13>.NET_003 0 0.183127f
c_97288 XI1.XI0.XI1<7>.XI7<13>.NET_005 0 0.0724835f
c_97307 XI1.XI0.XI1<7>.XI7<12>.NET_000 0 0.191272f
c_97322 XI1.XI0.XI1<7>.XI7<12>.NET_001 0 0.0667363f
c_97339 XI1.XI0.XI1<7>.XI7<12>.NET_003 0 0.184437f
c_97354 XI1.XI0.XI1<7>.XI7<12>.NET_005 0 0.0732094f
c_97376 XI1.XI0.XI1<6>.XI7<3>.NET_000 0 0.187391f
c_97394 XI1.XI0.XI1<6>.XI7<3>.NET_001 0 0.0680399f
c_97413 XI1.XI0.XI1<6>.XI7<3>.NET_003 0 0.181648f
c_97428 XI1.XI0.XI1<6>.XI7<3>.NET_005 0 0.0740537f
c_97449 XI1.XI0.XI1<6>.XI7<2>.NET_000 0 0.187429f
c_97467 XI1.XI0.XI1<6>.XI7<2>.NET_001 0 0.0670282f
c_97486 XI1.XI0.XI1<6>.XI7<2>.NET_003 0 0.180907f
c_97501 XI1.XI0.XI1<6>.XI7<2>.NET_005 0 0.0740537f
c_97523 XI1.XI0.XI1<6>.XI7<1>.NET_000 0 0.186614f
c_97541 XI1.XI0.XI1<6>.XI7<1>.NET_001 0 0.0675769f
c_97560 XI1.XI0.XI1<6>.XI7<1>.NET_003 0 0.181754f
c_97575 XI1.XI0.XI1<6>.XI7<1>.NET_005 0 0.0740537f
c_97597 XI1.XI0.XI1<6>.XI7<0>.NET_000 0 0.191342f
c_97614 XI1.XI0.XI1<6>.XI7<0>.NET_001 0 0.0672192f
c_97633 XI1.XI0.XI1<6>.XI7<0>.NET_003 0 0.18234f
c_97648 XI1.XI0.XI1<6>.XI7<0>.NET_005 0 0.0740681f
c_97667 XI1.XI0.XI1<6>.XI7<7>.NET_000 0 0.197638f
c_97684 XI1.XI0.XI1<6>.XI7<7>.NET_001 0 0.0680332f
c_97701 XI1.XI0.XI1<6>.XI7<7>.NET_003 0 0.18397f
c_97716 XI1.XI0.XI1<6>.XI7<7>.NET_005 0 0.0740187f
c_97735 XI1.XI0.XI1<6>.XI7<6>.NET_000 0 0.189436f
c_97751 XI1.XI0.XI1<6>.XI7<6>.NET_001 0 0.0671634f
c_97768 XI1.XI0.XI1<6>.XI7<6>.NET_003 0 0.181559f
c_97783 XI1.XI0.XI1<6>.XI7<6>.NET_005 0 0.0740537f
c_97804 XI1.XI0.XI1<6>.XI7<5>.NET_000 0 0.18932f
c_97821 XI1.XI0.XI1<6>.XI7<5>.NET_001 0 0.0678117f
c_97840 XI1.XI0.XI1<6>.XI7<5>.NET_003 0 0.182281f
c_97855 XI1.XI0.XI1<6>.XI7<5>.NET_005 0 0.0740537f
c_97875 XI1.XI0.XI1<6>.XI7<4>.NET_000 0 0.18791f
c_97891 XI1.XI0.XI1<6>.XI7<4>.NET_001 0 0.0676945f
c_97909 XI1.XI0.XI1<6>.XI7<4>.NET_003 0 0.180953f
c_97924 XI1.XI0.XI1<6>.XI7<4>.NET_005 0 0.0740537f
c_97943 XI1.XI0.XI1<6>.XI7<11>.NET_000 0 0.189304f
c_97958 XI1.XI0.XI1<6>.XI7<11>.NET_001 0 0.0685193f
c_97974 XI1.XI0.XI1<6>.XI7<11>.NET_003 0 0.182476f
c_97990 XI1.XI0.XI1<6>.XI7<11>.NET_005 0 0.0724229f
c_98009 XI1.XI0.XI1<6>.XI7<10>.NET_000 0 0.190142f
c_98024 XI1.XI0.XI1<6>.XI7<10>.NET_001 0 0.0671183f
c_98041 XI1.XI0.XI1<6>.XI7<10>.NET_003 0 0.182771f
c_98057 XI1.XI0.XI1<6>.XI7<10>.NET_005 0 0.0724229f
c_98077 XI1.XI0.XI1<6>.XI7<9>.NET_000 0 0.189836f
c_98093 XI1.XI0.XI1<6>.XI7<9>.NET_001 0 0.0683151f
c_98111 XI1.XI0.XI1<6>.XI7<9>.NET_003 0 0.182339f
c_98127 XI1.XI0.XI1<6>.XI7<9>.NET_005 0 0.0724229f
c_98149 XI1.XI0.XI1<6>.XI7<8>.NET_000 0 0.195684f
c_98165 XI1.XI0.XI1<6>.XI7<8>.NET_001 0 0.0669071f
c_98182 XI1.XI0.XI1<6>.XI7<8>.NET_003 0 0.181615f
c_98198 XI1.XI0.XI1<6>.XI7<8>.NET_005 0 0.0721499f
c_98218 XI1.XI0.XI1<6>.XI7<15>.NET_000 0 0.190105f
c_98235 XI1.XI0.XI1<6>.XI7<15>.NET_001 0 0.0677275f
c_98252 XI1.XI0.XI1<6>.XI7<15>.NET_003 0 0.182845f
c_98268 XI1.XI0.XI1<6>.XI7<15>.NET_005 0 0.0726863f
c_98290 XI1.XI0.XI1<6>.XI7<14>.NET_000 0 0.18727f
c_98308 XI1.XI0.XI1<6>.XI7<14>.NET_001 0 0.0669549f
c_98327 XI1.XI0.XI1<6>.XI7<14>.NET_003 0 0.181213f
c_98343 XI1.XI0.XI1<6>.XI7<14>.NET_005 0 0.0724229f
c_98363 XI1.XI0.XI1<6>.XI7<13>.NET_000 0 0.18825f
c_98379 XI1.XI0.XI1<6>.XI7<13>.NET_001 0 0.0689289f
c_98396 XI1.XI0.XI1<6>.XI7<13>.NET_003 0 0.183155f
c_98412 XI1.XI0.XI1<6>.XI7<13>.NET_005 0 0.0724623f
c_98432 XI1.XI0.XI1<6>.XI7<12>.NET_000 0 0.191236f
c_98448 XI1.XI0.XI1<6>.XI7<12>.NET_001 0 0.0667198f
c_98465 XI1.XI0.XI1<6>.XI7<12>.NET_003 0 0.184444f
c_98480 XI1.XI0.XI1<6>.XI7<12>.NET_005 0 0.0731882f
c_98502 XI1.XI0.XI1<5>.XI7<3>.NET_000 0 0.187617f
c_98520 XI1.XI0.XI1<5>.XI7<3>.NET_001 0 0.0680399f
c_98539 XI1.XI0.XI1<5>.XI7<3>.NET_003 0 0.18167f
c_98554 XI1.XI0.XI1<5>.XI7<3>.NET_005 0 0.0724441f
c_98575 XI1.XI0.XI1<5>.XI7<2>.NET_000 0 0.187648f
c_98593 XI1.XI0.XI1<5>.XI7<2>.NET_001 0 0.0670282f
c_98612 XI1.XI0.XI1<5>.XI7<2>.NET_003 0 0.180907f
c_98627 XI1.XI0.XI1<5>.XI7<2>.NET_005 0 0.0724441f
c_98649 XI1.XI0.XI1<5>.XI7<1>.NET_000 0 0.186864f
c_98667 XI1.XI0.XI1<5>.XI7<1>.NET_001 0 0.0676071f
c_98686 XI1.XI0.XI1<5>.XI7<1>.NET_003 0 0.181857f
c_98701 XI1.XI0.XI1<5>.XI7<1>.NET_005 0 0.0724441f
c_98722 XI1.XI0.XI1<5>.XI7<0>.NET_000 0 0.19148f
c_98738 XI1.XI0.XI1<5>.XI7<0>.NET_001 0 0.0672494f
c_98756 XI1.XI0.XI1<5>.XI7<0>.NET_003 0 0.182489f
c_98772 XI1.XI0.XI1<5>.XI7<0>.NET_005 0 0.0724585f
c_98791 XI1.XI0.XI1<5>.XI7<7>.NET_000 0 0.197939f
c_98808 XI1.XI0.XI1<5>.XI7<7>.NET_001 0 0.0679843f
c_98825 XI1.XI0.XI1<5>.XI7<7>.NET_003 0 0.183962f
c_98840 XI1.XI0.XI1<5>.XI7<7>.NET_005 0 0.0724512f
c_98859 XI1.XI0.XI1<5>.XI7<6>.NET_000 0 0.189655f
c_98875 XI1.XI0.XI1<5>.XI7<6>.NET_001 0 0.0671634f
c_98892 XI1.XI0.XI1<5>.XI7<6>.NET_003 0 0.181559f
c_98907 XI1.XI0.XI1<5>.XI7<6>.NET_005 0 0.0724441f
c_98928 XI1.XI0.XI1<5>.XI7<5>.NET_000 0 0.189539f
c_98945 XI1.XI0.XI1<5>.XI7<5>.NET_001 0 0.0678117f
c_98964 XI1.XI0.XI1<5>.XI7<5>.NET_003 0 0.182305f
c_98979 XI1.XI0.XI1<5>.XI7<5>.NET_005 0 0.0724441f
c_98999 XI1.XI0.XI1<5>.XI7<4>.NET_000 0 0.188128f
c_99015 XI1.XI0.XI1<5>.XI7<4>.NET_001 0 0.0676945f
c_99033 XI1.XI0.XI1<5>.XI7<4>.NET_003 0 0.180953f
c_99048 XI1.XI0.XI1<5>.XI7<4>.NET_005 0 0.0724441f
c_99066 XI1.XI0.XI1<5>.XI7<11>.NET_000 0 0.189523f
c_99081 XI1.XI0.XI1<5>.XI7<11>.NET_001 0 0.0685193f
c_99097 XI1.XI0.XI1<5>.XI7<11>.NET_003 0 0.182476f
c_99113 XI1.XI0.XI1<5>.XI7<11>.NET_005 0 0.0724441f
c_99132 XI1.XI0.XI1<5>.XI7<10>.NET_000 0 0.190324f
c_99148 XI1.XI0.XI1<5>.XI7<10>.NET_001 0 0.0671019f
c_99165 XI1.XI0.XI1<5>.XI7<10>.NET_003 0 0.182778f
c_99181 XI1.XI0.XI1<5>.XI7<10>.NET_005 0 0.0724441f
c_99200 XI1.XI0.XI1<5>.XI7<9>.NET_000 0 0.190054f
c_99216 XI1.XI0.XI1<5>.XI7<9>.NET_001 0 0.0683151f
c_99233 XI1.XI0.XI1<5>.XI7<9>.NET_003 0 0.182367f
c_99249 XI1.XI0.XI1<5>.XI7<9>.NET_005 0 0.0724441f
c_99270 XI1.XI0.XI1<5>.XI7<8>.NET_000 0 0.195902f
c_99286 XI1.XI0.XI1<5>.XI7<8>.NET_001 0 0.0669071f
c_99304 XI1.XI0.XI1<5>.XI7<8>.NET_003 0 0.181592f
c_99320 XI1.XI0.XI1<5>.XI7<8>.NET_005 0 0.0721711f
c_99339 XI1.XI0.XI1<5>.XI7<15>.NET_000 0 0.190352f
c_99356 XI1.XI0.XI1<5>.XI7<15>.NET_001 0 0.0677275f
c_99373 XI1.XI0.XI1<5>.XI7<15>.NET_003 0 0.182845f
c_99389 XI1.XI0.XI1<5>.XI7<15>.NET_005 0 0.0727082f
c_99410 XI1.XI0.XI1<5>.XI7<14>.NET_000 0 0.187509f
c_99428 XI1.XI0.XI1<5>.XI7<14>.NET_001 0 0.0669564f
c_99447 XI1.XI0.XI1<5>.XI7<14>.NET_003 0 0.181224f
c_99463 XI1.XI0.XI1<5>.XI7<14>.NET_005 0 0.0724441f
c_99482 XI1.XI0.XI1<5>.XI7<13>.NET_000 0 0.188468f
c_99498 XI1.XI0.XI1<5>.XI7<13>.NET_001 0 0.0689289f
c_99515 XI1.XI0.XI1<5>.XI7<13>.NET_003 0 0.183155f
c_99531 XI1.XI0.XI1<5>.XI7<13>.NET_005 0 0.0724835f
c_99550 XI1.XI0.XI1<5>.XI7<12>.NET_000 0 0.19145f
c_99566 XI1.XI0.XI1<5>.XI7<12>.NET_001 0 0.0667214f
c_99583 XI1.XI0.XI1<5>.XI7<12>.NET_003 0 0.184454f
c_99598 XI1.XI0.XI1<5>.XI7<12>.NET_005 0 0.0732094f
c_99620 XI1.XI0.XI1<4>.XI7<3>.NET_000 0 0.187398f
c_99638 XI1.XI0.XI1<4>.XI7<3>.NET_001 0 0.0680399f
c_99657 XI1.XI0.XI1<4>.XI7<3>.NET_003 0 0.181695f
c_99672 XI1.XI0.XI1<4>.XI7<3>.NET_005 0 0.0724441f
c_99693 XI1.XI0.XI1<4>.XI7<2>.NET_000 0 0.187429f
c_99711 XI1.XI0.XI1<4>.XI7<2>.NET_001 0 0.0670282f
c_99730 XI1.XI0.XI1<4>.XI7<2>.NET_003 0 0.180907f
c_99745 XI1.XI0.XI1<4>.XI7<2>.NET_005 0 0.0724441f
c_99767 XI1.XI0.XI1<4>.XI7<1>.NET_000 0 0.186653f
c_99785 XI1.XI0.XI1<4>.XI7<1>.NET_001 0 0.0676071f
c_99804 XI1.XI0.XI1<4>.XI7<1>.NET_003 0 0.181879f
c_99819 XI1.XI0.XI1<4>.XI7<1>.NET_005 0 0.0724441f
c_99840 XI1.XI0.XI1<4>.XI7<0>.NET_000 0 0.191381f
c_99856 XI1.XI0.XI1<4>.XI7<0>.NET_001 0 0.0672494f
c_99874 XI1.XI0.XI1<4>.XI7<0>.NET_003 0 0.182489f
c_99890 XI1.XI0.XI1<4>.XI7<0>.NET_005 0 0.0724585f
c_99909 XI1.XI0.XI1<4>.XI7<7>.NET_000 0 0.197616f
c_99926 XI1.XI0.XI1<4>.XI7<7>.NET_001 0 0.0679353f
c_99943 XI1.XI0.XI1<4>.XI7<7>.NET_003 0 0.183957f
c_99958 XI1.XI0.XI1<4>.XI7<7>.NET_005 0 0.0724512f
c_99977 XI1.XI0.XI1<4>.XI7<6>.NET_000 0 0.189436f
c_99993 XI1.XI0.XI1<4>.XI7<6>.NET_001 0 0.0671634f
c_100010 XI1.XI0.XI1<4>.XI7<6>.NET_003 0 0.181559f
c_100025 XI1.XI0.XI1<4>.XI7<6>.NET_005 0 0.0724441f
c_100046 XI1.XI0.XI1<4>.XI7<5>.NET_000 0 0.189304f
c_100063 XI1.XI0.XI1<4>.XI7<5>.NET_001 0 0.0678117f
c_100082 XI1.XI0.XI1<4>.XI7<5>.NET_003 0 0.182295f
c_100097 XI1.XI0.XI1<4>.XI7<5>.NET_005 0 0.0724441f
c_100117 XI1.XI0.XI1<4>.XI7<4>.NET_000 0 0.18791f
c_100133 XI1.XI0.XI1<4>.XI7<4>.NET_001 0 0.0676945f
c_100151 XI1.XI0.XI1<4>.XI7<4>.NET_003 0 0.180953f
c_100166 XI1.XI0.XI1<4>.XI7<4>.NET_005 0 0.0724441f
c_100185 XI1.XI0.XI1<4>.XI7<11>.NET_000 0 0.189304f
c_100200 XI1.XI0.XI1<4>.XI7<11>.NET_001 0 0.0685193f
c_100216 XI1.XI0.XI1<4>.XI7<11>.NET_003 0 0.182476f
c_100232 XI1.XI0.XI1<4>.XI7<11>.NET_005 0 0.0724441f
c_100252 XI1.XI0.XI1<4>.XI7<10>.NET_000 0 0.190126f
c_100268 XI1.XI0.XI1<4>.XI7<10>.NET_001 0 0.0671034f
c_100285 XI1.XI0.XI1<4>.XI7<10>.NET_003 0 0.182788f
c_100301 XI1.XI0.XI1<4>.XI7<10>.NET_005 0 0.0724441f
c_100321 XI1.XI0.XI1<4>.XI7<9>.NET_000 0 0.189836f
c_100337 XI1.XI0.XI1<4>.XI7<9>.NET_001 0 0.0683151f
c_100354 XI1.XI0.XI1<4>.XI7<9>.NET_003 0 0.182367f
c_100370 XI1.XI0.XI1<4>.XI7<9>.NET_005 0 0.0724441f
c_100393 XI1.XI0.XI1<4>.XI7<8>.NET_000 0 0.19558f
c_100410 XI1.XI0.XI1<4>.XI7<8>.NET_001 0 0.0668887f
c_100428 XI1.XI0.XI1<4>.XI7<8>.NET_003 0 0.181604f
c_100444 XI1.XI0.XI1<4>.XI7<8>.NET_005 0 0.0721711f
c_100464 XI1.XI0.XI1<4>.XI7<15>.NET_000 0 0.190105f
c_100481 XI1.XI0.XI1<4>.XI7<15>.NET_001 0 0.0677275f
c_100498 XI1.XI0.XI1<4>.XI7<15>.NET_003 0 0.182845f
c_100514 XI1.XI0.XI1<4>.XI7<15>.NET_005 0 0.0727082f
c_100536 XI1.XI0.XI1<4>.XI7<14>.NET_000 0 0.187306f
c_100554 XI1.XI0.XI1<4>.XI7<14>.NET_001 0 0.0669713f
c_100573 XI1.XI0.XI1<4>.XI7<14>.NET_003 0 0.18123f
c_100589 XI1.XI0.XI1<4>.XI7<14>.NET_005 0 0.0724441f
c_100609 XI1.XI0.XI1<4>.XI7<13>.NET_000 0 0.18825f
c_100625 XI1.XI0.XI1<4>.XI7<13>.NET_001 0 0.0689289f
c_100642 XI1.XI0.XI1<4>.XI7<13>.NET_003 0 0.183155f
c_100658 XI1.XI0.XI1<4>.XI7<13>.NET_005 0 0.0724835f
c_100678 XI1.XI0.XI1<4>.XI7<12>.NET_000 0 0.191272f
c_100694 XI1.XI0.XI1<4>.XI7<12>.NET_001 0 0.0667363f
c_100711 XI1.XI0.XI1<4>.XI7<12>.NET_003 0 0.184465f
c_100726 XI1.XI0.XI1<4>.XI7<12>.NET_005 0 0.0732094f
c_100748 XI1.XI0.XI1<3>.XI7<3>.NET_000 0 0.187383f
c_100766 XI1.XI0.XI1<3>.XI7<3>.NET_001 0 0.0680399f
c_100785 XI1.XI0.XI1<3>.XI7<3>.NET_003 0 0.181695f
c_100800 XI1.XI0.XI1<3>.XI7<3>.NET_005 0 0.0724441f
c_100821 XI1.XI0.XI1<3>.XI7<2>.NET_000 0 0.187429f
c_100839 XI1.XI0.XI1<3>.XI7<2>.NET_001 0 0.0670282f
c_100858 XI1.XI0.XI1<3>.XI7<2>.NET_003 0 0.180907f
c_100873 XI1.XI0.XI1<3>.XI7<2>.NET_005 0 0.0724441f
c_100895 XI1.XI0.XI1<3>.XI7<1>.NET_000 0 0.186653f
c_100913 XI1.XI0.XI1<3>.XI7<1>.NET_001 0 0.0676071f
c_100932 XI1.XI0.XI1<3>.XI7<1>.NET_003 0 0.181903f
c_100947 XI1.XI0.XI1<3>.XI7<1>.NET_005 0 0.0724441f
c_100968 XI1.XI0.XI1<3>.XI7<0>.NET_000 0 0.191381f
c_100984 XI1.XI0.XI1<3>.XI7<0>.NET_001 0 0.0672494f
c_101002 XI1.XI0.XI1<3>.XI7<0>.NET_003 0 0.182489f
c_101018 XI1.XI0.XI1<3>.XI7<0>.NET_005 0 0.0724585f
c_101036 XI1.XI0.XI1<3>.XI7<7>.NET_000 0 0.197811f
c_101052 XI1.XI0.XI1<3>.XI7<7>.NET_001 0 0.0680452f
c_101069 XI1.XI0.XI1<3>.XI7<7>.NET_003 0 0.183961f
c_101084 XI1.XI0.XI1<3>.XI7<7>.NET_005 0 0.0724146f
c_101103 XI1.XI0.XI1<3>.XI7<6>.NET_000 0 0.189436f
c_101119 XI1.XI0.XI1<3>.XI7<6>.NET_001 0 0.0671634f
c_101136 XI1.XI0.XI1<3>.XI7<6>.NET_003 0 0.181559f
c_101151 XI1.XI0.XI1<3>.XI7<6>.NET_005 0 0.0724441f
c_101172 XI1.XI0.XI1<3>.XI7<5>.NET_000 0 0.189284f
c_101189 XI1.XI0.XI1<3>.XI7<5>.NET_001 0 0.0678117f
c_101208 XI1.XI0.XI1<3>.XI7<5>.NET_003 0 0.182284f
c_101223 XI1.XI0.XI1<3>.XI7<5>.NET_005 0 0.0724441f
c_101243 XI1.XI0.XI1<3>.XI7<4>.NET_000 0 0.18791f
c_101259 XI1.XI0.XI1<3>.XI7<4>.NET_001 0 0.0676945f
c_101277 XI1.XI0.XI1<3>.XI7<4>.NET_003 0 0.180953f
c_101292 XI1.XI0.XI1<3>.XI7<4>.NET_005 0 0.0724441f
c_101311 XI1.XI0.XI1<3>.XI7<11>.NET_000 0 0.189304f
c_101326 XI1.XI0.XI1<3>.XI7<11>.NET_001 0 0.0685193f
c_101342 XI1.XI0.XI1<3>.XI7<11>.NET_003 0 0.182476f
c_101358 XI1.XI0.XI1<3>.XI7<11>.NET_005 0 0.0724441f
c_101378 XI1.XI0.XI1<3>.XI7<10>.NET_000 0 0.190142f
c_101394 XI1.XI0.XI1<3>.XI7<10>.NET_001 0 0.0671183f
c_101411 XI1.XI0.XI1<3>.XI7<10>.NET_003 0 0.182799f
c_101427 XI1.XI0.XI1<3>.XI7<10>.NET_005 0 0.0724441f
c_101447 XI1.XI0.XI1<3>.XI7<9>.NET_000 0 0.189836f
c_101463 XI1.XI0.XI1<3>.XI7<9>.NET_001 0 0.0683151f
c_101480 XI1.XI0.XI1<3>.XI7<9>.NET_003 0 0.182367f
c_101496 XI1.XI0.XI1<3>.XI7<9>.NET_005 0 0.0724441f
c_101519 XI1.XI0.XI1<3>.XI7<8>.NET_000 0 0.195684f
c_101536 XI1.XI0.XI1<3>.XI7<8>.NET_001 0 0.0669071f
c_101554 XI1.XI0.XI1<3>.XI7<8>.NET_003 0 0.181619f
c_101570 XI1.XI0.XI1<3>.XI7<8>.NET_005 0 0.0721711f
c_101590 XI1.XI0.XI1<3>.XI7<15>.NET_000 0 0.190105f
c_101607 XI1.XI0.XI1<3>.XI7<15>.NET_001 0 0.0677275f
c_101624 XI1.XI0.XI1<3>.XI7<15>.NET_003 0 0.182845f
c_101640 XI1.XI0.XI1<3>.XI7<15>.NET_005 0 0.0727082f
c_101662 XI1.XI0.XI1<3>.XI7<14>.NET_000 0 0.187306f
c_101680 XI1.XI0.XI1<3>.XI7<14>.NET_001 0 0.0669713f
c_101699 XI1.XI0.XI1<3>.XI7<14>.NET_003 0 0.18121f
c_101715 XI1.XI0.XI1<3>.XI7<14>.NET_005 0 0.0724441f
c_101735 XI1.XI0.XI1<3>.XI7<13>.NET_000 0 0.18825f
c_101751 XI1.XI0.XI1<3>.XI7<13>.NET_001 0 0.0689289f
c_101768 XI1.XI0.XI1<3>.XI7<13>.NET_003 0 0.183155f
c_101784 XI1.XI0.XI1<3>.XI7<13>.NET_005 0 0.0724835f
c_101804 XI1.XI0.XI1<3>.XI7<12>.NET_000 0 0.191272f
c_101820 XI1.XI0.XI1<3>.XI7<12>.NET_001 0 0.0667363f
c_101837 XI1.XI0.XI1<3>.XI7<12>.NET_003 0 0.18446f
c_101852 XI1.XI0.XI1<3>.XI7<12>.NET_005 0 0.0732094f
c_101874 XI1.XI0.XI1<2>.XI7<3>.NET_000 0 0.187362f
c_101892 XI1.XI0.XI1<2>.XI7<3>.NET_001 0 0.0680399f
c_101911 XI1.XI0.XI1<2>.XI7<3>.NET_003 0 0.181695f
c_101926 XI1.XI0.XI1<2>.XI7<3>.NET_005 0 0.0724441f
c_101947 XI1.XI0.XI1<2>.XI7<2>.NET_000 0 0.187429f
c_101965 XI1.XI0.XI1<2>.XI7<2>.NET_001 0 0.0670282f
c_101984 XI1.XI0.XI1<2>.XI7<2>.NET_003 0 0.180907f
c_101999 XI1.XI0.XI1<2>.XI7<2>.NET_005 0 0.0724441f
c_102021 XI1.XI0.XI1<2>.XI7<1>.NET_000 0 0.186653f
c_102039 XI1.XI0.XI1<2>.XI7<1>.NET_001 0 0.0676071f
c_102058 XI1.XI0.XI1<2>.XI7<1>.NET_003 0 0.181903f
c_102073 XI1.XI0.XI1<2>.XI7<1>.NET_005 0 0.0724441f
c_102094 XI1.XI0.XI1<2>.XI7<0>.NET_000 0 0.191381f
c_102110 XI1.XI0.XI1<2>.XI7<0>.NET_001 0 0.0672494f
c_102128 XI1.XI0.XI1<2>.XI7<0>.NET_003 0 0.182489f
c_102144 XI1.XI0.XI1<2>.XI7<0>.NET_005 0 0.0724585f
c_102162 XI1.XI0.XI1<2>.XI7<7>.NET_000 0 0.197681f
c_102178 XI1.XI0.XI1<2>.XI7<7>.NET_001 0 0.0680197f
c_102194 XI1.XI0.XI1<2>.XI7<7>.NET_003 0 0.183965f
c_102209 XI1.XI0.XI1<2>.XI7<7>.NET_005 0 0.0724585f
c_102228 XI1.XI0.XI1<2>.XI7<6>.NET_000 0 0.189436f
c_102244 XI1.XI0.XI1<2>.XI7<6>.NET_001 0 0.0671634f
c_102262 XI1.XI0.XI1<2>.XI7<6>.NET_003 0 0.181531f
c_102277 XI1.XI0.XI1<2>.XI7<6>.NET_005 0 0.0724441f
c_102297 XI1.XI0.XI1<2>.XI7<5>.NET_000 0 0.18932f
c_102314 XI1.XI0.XI1<2>.XI7<5>.NET_001 0 0.0678117f
c_102333 XI1.XI0.XI1<2>.XI7<5>.NET_003 0 0.182278f
c_102348 XI1.XI0.XI1<2>.XI7<5>.NET_005 0 0.0724441f
c_102368 XI1.XI0.XI1<2>.XI7<4>.NET_000 0 0.18791f
c_102384 XI1.XI0.XI1<2>.XI7<4>.NET_001 0 0.0676945f
c_102402 XI1.XI0.XI1<2>.XI7<4>.NET_003 0 0.180953f
c_102417 XI1.XI0.XI1<2>.XI7<4>.NET_005 0 0.0724441f
c_102436 XI1.XI0.XI1<2>.XI7<11>.NET_000 0 0.189304f
c_102451 XI1.XI0.XI1<2>.XI7<11>.NET_001 0 0.0685193f
c_102467 XI1.XI0.XI1<2>.XI7<11>.NET_003 0 0.182476f
c_102483 XI1.XI0.XI1<2>.XI7<11>.NET_005 0 0.0724441f
c_102503 XI1.XI0.XI1<2>.XI7<10>.NET_000 0 0.190142f
c_102519 XI1.XI0.XI1<2>.XI7<10>.NET_001 0 0.0671183f
c_102536 XI1.XI0.XI1<2>.XI7<10>.NET_003 0 0.182799f
c_102552 XI1.XI0.XI1<2>.XI7<10>.NET_005 0 0.0724441f
c_102572 XI1.XI0.XI1<2>.XI7<9>.NET_000 0 0.189836f
c_102588 XI1.XI0.XI1<2>.XI7<9>.NET_001 0 0.0683151f
c_102605 XI1.XI0.XI1<2>.XI7<9>.NET_003 0 0.182367f
c_102621 XI1.XI0.XI1<2>.XI7<9>.NET_005 0 0.0724441f
c_102644 XI1.XI0.XI1<2>.XI7<8>.NET_000 0 0.195684f
c_102661 XI1.XI0.XI1<2>.XI7<8>.NET_001 0 0.0669071f
c_102679 XI1.XI0.XI1<2>.XI7<8>.NET_003 0 0.181619f
c_102695 XI1.XI0.XI1<2>.XI7<8>.NET_005 0 0.0721711f
c_102715 XI1.XI0.XI1<2>.XI7<15>.NET_000 0 0.190105f
c_102732 XI1.XI0.XI1<2>.XI7<15>.NET_001 0 0.0677275f
c_102749 XI1.XI0.XI1<2>.XI7<15>.NET_003 0 0.182845f
c_102765 XI1.XI0.XI1<2>.XI7<15>.NET_005 0 0.0727082f
c_102787 XI1.XI0.XI1<2>.XI7<14>.NET_000 0 0.187299f
c_102805 XI1.XI0.XI1<2>.XI7<14>.NET_001 0 0.0669713f
c_102824 XI1.XI0.XI1<2>.XI7<14>.NET_003 0 0.181188f
c_102840 XI1.XI0.XI1<2>.XI7<14>.NET_005 0 0.0724441f
c_102860 XI1.XI0.XI1<2>.XI7<13>.NET_000 0 0.18825f
c_102876 XI1.XI0.XI1<2>.XI7<13>.NET_001 0 0.0689289f
c_102893 XI1.XI0.XI1<2>.XI7<13>.NET_003 0 0.183155f
c_102909 XI1.XI0.XI1<2>.XI7<13>.NET_005 0 0.0724835f
c_102929 XI1.XI0.XI1<2>.XI7<12>.NET_000 0 0.191272f
c_102945 XI1.XI0.XI1<2>.XI7<12>.NET_001 0 0.0667363f
c_102962 XI1.XI0.XI1<2>.XI7<12>.NET_003 0 0.18444f
c_102977 XI1.XI0.XI1<2>.XI7<12>.NET_005 0 0.0732094f
c_102998 XI1.XI0.XI1<1>.XI7<3>.NET_000 0 0.187398f
c_103016 XI1.XI0.XI1<1>.XI7<3>.NET_001 0 0.0680399f
c_103035 XI1.XI0.XI1<1>.XI7<3>.NET_003 0 0.181695f
c_103050 XI1.XI0.XI1<1>.XI7<3>.NET_005 0 0.0724441f
c_103071 XI1.XI0.XI1<1>.XI7<2>.NET_000 0 0.187429f
c_103089 XI1.XI0.XI1<1>.XI7<2>.NET_001 0 0.0670282f
c_103108 XI1.XI0.XI1<1>.XI7<2>.NET_003 0 0.180907f
c_103123 XI1.XI0.XI1<1>.XI7<2>.NET_005 0 0.0724441f
c_103145 XI1.XI0.XI1<1>.XI7<1>.NET_000 0 0.186653f
c_103163 XI1.XI0.XI1<1>.XI7<1>.NET_001 0 0.0676071f
c_103182 XI1.XI0.XI1<1>.XI7<1>.NET_003 0 0.181903f
c_103197 XI1.XI0.XI1<1>.XI7<1>.NET_005 0 0.0724441f
c_103218 XI1.XI0.XI1<1>.XI7<0>.NET_000 0 0.191381f
c_103234 XI1.XI0.XI1<1>.XI7<0>.NET_001 0 0.0672494f
c_103252 XI1.XI0.XI1<1>.XI7<0>.NET_003 0 0.182489f
c_103268 XI1.XI0.XI1<1>.XI7<0>.NET_005 0 0.0724585f
c_103286 XI1.XI0.XI1<1>.XI7<7>.NET_000 0 0.197741f
c_103302 XI1.XI0.XI1<1>.XI7<7>.NET_001 0 0.0680432f
c_103318 XI1.XI0.XI1<1>.XI7<7>.NET_003 0 0.184003f
c_103333 XI1.XI0.XI1<1>.XI7<7>.NET_005 0 0.0723985f
c_103353 XI1.XI0.XI1<1>.XI7<6>.NET_000 0 0.1894f
c_103370 XI1.XI0.XI1<1>.XI7<6>.NET_001 0 0.067147f
c_103388 XI1.XI0.XI1<1>.XI7<6>.NET_003 0 0.181538f
c_103403 XI1.XI0.XI1<1>.XI7<6>.NET_005 0 0.0724441f
c_103423 XI1.XI0.XI1<1>.XI7<5>.NET_000 0 0.18932f
c_103440 XI1.XI0.XI1<1>.XI7<5>.NET_001 0 0.0678117f
c_103458 XI1.XI0.XI1<1>.XI7<5>.NET_003 0 0.182305f
c_103473 XI1.XI0.XI1<1>.XI7<5>.NET_005 0 0.0724441f
c_103493 XI1.XI0.XI1<1>.XI7<4>.NET_000 0 0.18791f
c_103509 XI1.XI0.XI1<1>.XI7<4>.NET_001 0 0.0676945f
c_103528 XI1.XI0.XI1<1>.XI7<4>.NET_003 0 0.180925f
c_103543 XI1.XI0.XI1<1>.XI7<4>.NET_005 0 0.0724441f
c_103562 XI1.XI0.XI1<1>.XI7<11>.NET_000 0 0.189304f
c_103577 XI1.XI0.XI1<1>.XI7<11>.NET_001 0 0.0685193f
c_103593 XI1.XI0.XI1<1>.XI7<11>.NET_003 0 0.182476f
c_103609 XI1.XI0.XI1<1>.XI7<11>.NET_005 0 0.0724441f
c_103629 XI1.XI0.XI1<1>.XI7<10>.NET_000 0 0.190142f
c_103645 XI1.XI0.XI1<1>.XI7<10>.NET_001 0 0.0671183f
c_103662 XI1.XI0.XI1<1>.XI7<10>.NET_003 0 0.182799f
c_103678 XI1.XI0.XI1<1>.XI7<10>.NET_005 0 0.0724441f
c_103698 XI1.XI0.XI1<1>.XI7<9>.NET_000 0 0.189836f
c_103714 XI1.XI0.XI1<1>.XI7<9>.NET_001 0 0.0683151f
c_103731 XI1.XI0.XI1<1>.XI7<9>.NET_003 0 0.182367f
c_103747 XI1.XI0.XI1<1>.XI7<9>.NET_005 0 0.0724441f
c_103770 XI1.XI0.XI1<1>.XI7<8>.NET_000 0 0.195684f
c_103787 XI1.XI0.XI1<1>.XI7<8>.NET_001 0 0.0669071f
c_103805 XI1.XI0.XI1<1>.XI7<8>.NET_003 0 0.181619f
c_103821 XI1.XI0.XI1<1>.XI7<8>.NET_005 0 0.0721711f
c_103842 XI1.XI0.XI1<1>.XI7<15>.NET_000 0 0.190066f
c_103860 XI1.XI0.XI1<1>.XI7<15>.NET_001 0 0.0676964f
c_103878 XI1.XI0.XI1<1>.XI7<15>.NET_003 0 0.182696f
c_103894 XI1.XI0.XI1<1>.XI7<15>.NET_005 0 0.0727082f
c_103916 XI1.XI0.XI1<1>.XI7<14>.NET_000 0 0.187267f
c_103934 XI1.XI0.XI1<1>.XI7<14>.NET_001 0 0.0669403f
c_103953 XI1.XI0.XI1<1>.XI7<14>.NET_003 0 0.181085f
c_103969 XI1.XI0.XI1<1>.XI7<14>.NET_005 0 0.0724441f
c_103989 XI1.XI0.XI1<1>.XI7<13>.NET_000 0 0.18825f
c_104005 XI1.XI0.XI1<1>.XI7<13>.NET_001 0 0.0689289f
c_104022 XI1.XI0.XI1<1>.XI7<13>.NET_003 0 0.183155f
c_104038 XI1.XI0.XI1<1>.XI7<13>.NET_005 0 0.0724835f
c_104058 XI1.XI0.XI1<1>.XI7<12>.NET_000 0 0.191266f
c_104074 XI1.XI0.XI1<1>.XI7<12>.NET_001 0 0.0667363f
c_104091 XI1.XI0.XI1<1>.XI7<12>.NET_003 0 0.184419f
c_104106 XI1.XI0.XI1<1>.XI7<12>.NET_005 0 0.0732094f
c_104127 XI1.XI0.XI1<0>.XI7<3>.NET_000 0 0.187398f
c_104145 XI1.XI0.XI1<0>.XI7<3>.NET_001 0 0.0680945f
c_104164 XI1.XI0.XI1<0>.XI7<3>.NET_003 0 0.185169f
c_104180 XI1.XI0.XI1<0>.XI7<3>.NET_005 0 0.0776206f
c_104201 XI1.XI0.XI1<0>.XI7<2>.NET_000 0 0.187527f
c_104219 XI1.XI0.XI1<0>.XI7<2>.NET_001 0 0.0670356f
c_104239 XI1.XI0.XI1<0>.XI7<2>.NET_003 0 0.183267f
c_104253 XI1.XI0.XI1<0>.XI7<2>.NET_005 0 0.076804f
c_104275 XI1.XI0.XI1<0>.XI7<1>.NET_000 0 0.186653f
c_104293 XI1.XI0.XI1<0>.XI7<1>.NET_001 0 0.0676617f
c_104312 XI1.XI0.XI1<0>.XI7<1>.NET_003 0 0.185383f
c_104326 XI1.XI0.XI1<0>.XI7<1>.NET_005 0 0.0776206f
c_104347 XI1.XI0.XI1<0>.XI7<0>.NET_000 0 0.190934f
c_104363 XI1.XI0.XI1<0>.XI7<0>.NET_001 0 0.0672568f
c_104381 XI1.XI0.XI1<0>.XI7<0>.NET_003 0 0.184877f
c_104395 XI1.XI0.XI1<0>.XI7<0>.NET_005 0 0.0768185f
c_104413 XI1.XI0.XI1<0>.XI7<7>.NET_000 0 0.197619f
c_104429 XI1.XI0.XI1<0>.XI7<7>.NET_001 0 0.0678447f
c_104445 XI1.XI0.XI1<0>.XI7<7>.NET_003 0 0.187441f
c_104459 XI1.XI0.XI1<0>.XI7<7>.NET_005 0 0.0775644f
c_104479 XI1.XI0.XI1<0>.XI7<6>.NET_000 0 0.189519f
c_104496 XI1.XI0.XI1<0>.XI7<6>.NET_001 0 0.0671559f
c_104514 XI1.XI0.XI1<0>.XI7<6>.NET_003 0 0.183936f
c_104530 XI1.XI0.XI1<0>.XI7<6>.NET_005 0 0.076804f
c_104550 XI1.XI0.XI1<0>.XI7<5>.NET_000 0 0.18932f
c_104567 XI1.XI0.XI1<0>.XI7<5>.NET_001 0 0.0678663f
c_104585 XI1.XI0.XI1<0>.XI7<5>.NET_003 0 0.185785f
c_104602 XI1.XI0.XI1<0>.XI7<5>.NET_005 0 0.074256f
c_104623 XI1.XI0.XI1<0>.XI7<4>.NET_000 0 0.187972f
c_104640 XI1.XI0.XI1<0>.XI7<4>.NET_001 0 0.0676855f
c_104659 XI1.XI0.XI1<0>.XI7<4>.NET_003 0 0.18332f
c_104676 XI1.XI0.XI1<0>.XI7<4>.NET_005 0 0.0736665f
c_104696 XI1.XI0.XI1<0>.XI7<11>.NET_000 0 0.189265f
c_104712 XI1.XI0.XI1<0>.XI7<11>.NET_001 0 0.0685446f
c_104729 XI1.XI0.XI1<0>.XI7<11>.NET_003 0 0.185807f
c_104744 XI1.XI0.XI1<0>.XI7<11>.NET_005 0 0.0776206f
c_104764 XI1.XI0.XI1<0>.XI7<10>.NET_000 0 0.19024f
c_104780 XI1.XI0.XI1<0>.XI7<10>.NET_001 0 0.0671257f
c_104797 XI1.XI0.XI1<0>.XI7<10>.NET_003 0 0.185186f
c_104812 XI1.XI0.XI1<0>.XI7<10>.NET_005 0 0.076804f
c_104832 XI1.XI0.XI1<0>.XI7<9>.NET_000 0 0.189836f
c_104848 XI1.XI0.XI1<0>.XI7<9>.NET_001 0 0.0683696f
c_104865 XI1.XI0.XI1<0>.XI7<9>.NET_003 0 0.185847f
c_104880 XI1.XI0.XI1<0>.XI7<9>.NET_005 0 0.0776206f
c_104903 XI1.XI0.XI1<0>.XI7<8>.NET_000 0 0.195782f
c_104920 XI1.XI0.XI1<0>.XI7<8>.NET_001 0 0.0669268f
c_104938 XI1.XI0.XI1<0>.XI7<8>.NET_003 0 0.183997f
c_104953 XI1.XI0.XI1<0>.XI7<8>.NET_005 0 0.076531f
c_104974 XI1.XI0.XI1<0>.XI7<15>.NET_000 0 0.190087f
c_104992 XI1.XI0.XI1<0>.XI7<15>.NET_001 0 0.0677715f
c_105010 XI1.XI0.XI1<0>.XI7<15>.NET_003 0 0.186297f
c_105025 XI1.XI0.XI1<0>.XI7<15>.NET_005 0 0.077983f
c_105046 XI1.XI0.XI1<0>.XI7<14>.NET_000 0 0.187404f
c_105063 XI1.XI0.XI1<0>.XI7<14>.NET_001 0 0.0669787f
c_105081 XI1.XI0.XI1<0>.XI7<14>.NET_003 0 0.183622f
c_105098 XI1.XI0.XI1<0>.XI7<14>.NET_005 0 0.0767771f
c_105119 XI1.XI0.XI1<0>.XI7<13>.NET_000 0 0.18821f
c_105136 XI1.XI0.XI1<0>.XI7<13>.NET_001 0 0.0689541f
c_105154 XI1.XI0.XI1<0>.XI7<13>.NET_003 0 0.186485f
c_105172 XI1.XI0.XI1<0>.XI7<13>.NET_005 0 0.07766f
c_105192 XI1.XI0.XI1<0>.XI7<12>.NET_000 0 0.191331f
c_105208 XI1.XI0.XI1<0>.XI7<12>.NET_001 0 0.066724f
c_105225 XI1.XI0.XI1<0>.XI7<12>.NET_003 0 0.186797f
c_105239 XI1.XI0.XI1<0>.XI7<12>.NET_005 0 0.0775693f
c_105255 XI1.XI0.XI0.XI7<3>.NET_001 0 0.0822596f
c_105271 XI1.XI0.XI0.XI7<3>.NET_003 0 0.141475f
c_105285 XI1.XI0.XI0.XI7<3>.NET_005 0 0.055562f
c_105305 XI1.XI0.XI0.XI7<3>.NET_000 0 0.209745f
c_105321 XI1.XI0.XI0.XI7<2>.NET_001 0 0.0824899f
c_105337 XI1.XI0.XI0.XI7<2>.NET_003 0 0.142163f
c_105351 XI1.XI0.XI0.XI7<2>.NET_005 0 0.0557598f
c_105371 XI1.XI0.XI0.XI7<2>.NET_000 0 0.209746f
c_105387 XI1.XI0.XI0.XI7<1>.NET_001 0 0.0822596f
c_105403 XI1.XI0.XI0.XI7<1>.NET_003 0 0.141475f
c_105417 XI1.XI0.XI0.XI7<1>.NET_005 0 0.055562f
c_105437 XI1.XI0.XI0.XI7<1>.NET_000 0 0.209745f
c_105454 XI1.XI0.XI0.XI7<0>.NET_001 0 0.0825459f
c_105469 XI1.XI0.XI0.XI7<0>.NET_003 0 0.143041f
c_105483 XI1.XI0.XI0.XI7<0>.NET_005 0 0.0557446f
c_105503 XI1.XI0.XI0.XI7<0>.NET_000 0 0.222184f
c_105519 XI1.XI0.XI0.XI7<7>.NET_001 0 0.0823199f
c_105534 XI1.XI0.XI0.XI7<7>.NET_003 0 0.14235f
c_105548 XI1.XI0.XI0.XI7<7>.NET_005 0 0.0555395f
c_105568 XI1.XI0.XI0.XI7<7>.NET_000 0 0.222266f
c_105584 XI1.XI0.XI0.XI7<6>.NET_001 0 0.0824899f
c_105600 XI1.XI0.XI0.XI7<6>.NET_003 0 0.142163f
c_105614 XI1.XI0.XI0.XI7<6>.NET_005 0 0.0557598f
c_105634 XI1.XI0.XI0.XI7<6>.NET_000 0 0.209746f
c_105650 XI1.XI0.XI0.XI7<5>.NET_001 0 0.0822596f
c_105666 XI1.XI0.XI0.XI7<5>.NET_003 0 0.141475f
c_105680 XI1.XI0.XI0.XI7<5>.NET_005 0 0.055562f
c_105700 XI1.XI0.XI0.XI7<5>.NET_000 0 0.209745f
c_105716 XI1.XI0.XI0.XI7<4>.NET_001 0 0.0824899f
c_105732 XI1.XI0.XI0.XI7<4>.NET_003 0 0.142163f
c_105746 XI1.XI0.XI0.XI7<4>.NET_005 0 0.0557598f
c_105766 XI1.XI0.XI0.XI7<4>.NET_000 0 0.209746f
c_105782 XI1.XI0.XI0.XI7<11>.NET_001 0 0.0822596f
c_105798 XI1.XI0.XI0.XI7<11>.NET_003 0 0.141475f
c_105812 XI1.XI0.XI0.XI7<11>.NET_005 0 0.055562f
c_105833 XI1.XI0.XI0.XI7<11>.NET_000 0 0.209745f
c_105849 XI1.XI0.XI0.XI7<10>.NET_001 0 0.0824899f
c_105865 XI1.XI0.XI0.XI7<10>.NET_003 0 0.142163f
c_105879 XI1.XI0.XI0.XI7<10>.NET_005 0 0.0557598f
c_105900 XI1.XI0.XI0.XI7<10>.NET_000 0 0.209746f
c_105916 XI1.XI0.XI0.XI7<9>.NET_001 0 0.0822596f
c_105932 XI1.XI0.XI0.XI7<9>.NET_003 0 0.141475f
c_105946 XI1.XI0.XI0.XI7<9>.NET_005 0 0.055562f
c_105967 XI1.XI0.XI0.XI7<9>.NET_000 0 0.209745f
c_105983 XI1.XI0.XI0.XI7<8>.NET_001 0 0.08255f
c_105999 XI1.XI0.XI0.XI7<8>.NET_003 0 0.142643f
c_106013 XI1.XI0.XI0.XI7<8>.NET_005 0 0.0557622f
c_106040 XI1.XI0.XI0.XI7<8>.NET_000 0 0.219413f
c_106056 XI1.XI0.XI0.XI7<15>.NET_001 0 0.0826428f
c_106071 XI1.XI0.XI0.XI7<15>.NET_003 0 0.1422f
c_106084 XI1.XI0.XI0.XI7<15>.NET_005 0 0.0556175f
c_106105 XI1.XI0.XI0.XI7<15>.NET_000 0 0.222533f
c_106121 XI1.XI0.XI0.XI7<14>.NET_001 0 0.0824899f
c_106137 XI1.XI0.XI0.XI7<14>.NET_003 0 0.142163f
c_106151 XI1.XI0.XI0.XI7<14>.NET_005 0 0.0557598f
c_106172 XI1.XI0.XI0.XI7<14>.NET_000 0 0.209746f
c_106188 XI1.XI0.XI0.XI7<13>.NET_001 0 0.0822596f
c_106204 XI1.XI0.XI0.XI7<13>.NET_003 0 0.141569f
c_106218 XI1.XI0.XI0.XI7<13>.NET_005 0 0.055562f
c_106239 XI1.XI0.XI0.XI7<13>.NET_000 0 0.209745f
c_106254 XI1.XI0.XI0.XI7<12>.NET_001 0 0.0835715f
c_106269 XI1.XI0.XI0.XI7<12>.NET_003 0 0.144104f
c_106282 XI1.XI0.XI0.XI7<12>.NET_005 0 0.0565681f
c_106302 XI1.XI0.XI0.XI7<12>.NET_000 0 0.211123f
c_106313 XI1.XI0.XI21<1>.Z_NEG 0 0.148681f
c_106326 XI1.XI0.XI21<0>.Z_NEG 0 0.136548f
c_106341 XI1.XI0.XI20.Z_NEG 0 0.134909f
*
.include "RF.pex.netlist.RF.pxi"
*
.ends
*
*
