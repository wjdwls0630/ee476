* File: loaded_nand.pex.netlist
* Created: Fri Oct 29 05:31:21 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2
.subckt loaded_nand A B Z 
* 
mXDUT.MNMOS0 XDUT.NET2 A VSS! VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXDUT.MNMOS1 Z B XDUT.NET2 VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14
+ AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXDUT.MPMOS0 Z A VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14
+ PD=1.02e-06 PS=9.1e-07
mXDUT.MPMOS1 Z B VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14
+ PD=1.02e-06 PS=9.1e-07
mXI3.MNMOS0 XI3.NET2 VDD! VSS! VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI3.MNMOS1 NET4 Z XI3.NET2 VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14
+ AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXI3.MPMOS0 NET4 VDD! VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI3.MPMOS1 NET4 Z VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14
+ PD=1.02e-06 PS=9.1e-07
mXI2.MNMOS0 XI2.NET2 VDD! VSS! VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI2.MNMOS1 NET3 Z XI2.NET2 VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14
+ AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXI2.MPMOS0 NET3 VDD! VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI2.MPMOS1 NET3 Z VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14
+ PD=1.02e-06 PS=9.1e-07
mXI0.MNMOS0 XI0.NET2 VDD! VSS! VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI0.MNMOS1 NET2 Z XI0.NET2 VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14
+ AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXI0.MPMOS0 NET2 VDD! VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI0.MPMOS1 NET2 Z VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14
+ PD=1.02e-06 PS=9.1e-07
mXI1.MNMOS0 XI1.NET2 VDD! VSS! VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI1.MNMOS1 NET1 Z XI1.NET2 VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14
+ AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXI1.MPMOS0 NET1 VDD! VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI1.MPMOS1 NET1 Z VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14
+ PD=1.02e-06 PS=9.1e-07
c_9 Z 0 0.439259f
c_18 VDD! 0 0.866076f
c_23 A 0 0.0666759f
c_28 B 0 0.0637911f
c_37 VSS! 0 0.235132f
c_42 NET4 0 0.0196908f
c_47 NET3 0 0.0193199f
c_52 NET2 0 0.022558f
c_57 NET1 0 0.022558f
*
.include "loaded_nand.pex.netlist.LOADED_NAND.pxi"
*
.ends
*
*
