.GLOBAL vdd! vss!


.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2

* File: DFSR.pex.netlist
* Created: Mon Nov  8 16:45:41 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.include "DFSR.pex.netlist.pex"
.subckt DFSR CLK D Q RST 
* 
* CLK	CLK
* Q	Q
* D	D
* VSS!	VSS!
* VDD!	VDD!
* RST	RST
mXml0.Xnand0.MNMOS1 XML0.XNAND0.NET2 N_N_Xml0.Xnand0.MNMOS1_g
+ N_VSS!_Xml0.Xnand0.MNMOS1_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=2.5e-07
+ AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXml0.Xnand0.MNMOS0 N_XML0.N4_Xml0.Xnand0.MNMOS0_d
+ N_RST_BAR_Xml0.Xnand0.MNMOS0_g XML0.XNAND0.NET2 N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXsl0.Xnor0.MNMOS1 N_XSL0.N3_Xsl0.Xnor0.MNMOS1_d N_XSL0.N2_Xsl0.Xnor0.MNMOS1_g
+ N_VSS!_Xsl0.Xnor0.MNMOS1_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=9.5e-08
+ AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXsl0.Xnor0.MNMOS0 N_XSL0.N3_Xsl0.Xnor0.MNMOS1_d N_RST_Xsl0.Xnor0.MNMOS0_g
+ N_VSS!_Xsl0.Xnor0.MNMOS0_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=9.5e-08
+ AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXml0.Xnand0.MPMOS1 N_XML0.N4_Xml0.Xnand0.MPMOS1_d N_N_Xml0.Xnand0.MPMOS1_g
+ N_VDD!_Xml0.Xnand0.MPMOS1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=5.25e-07
+ AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXml0.Xnand0.MPMOS0 N_XML0.N4_Xml0.Xnand0.MPMOS1_d
+ N_RST_BAR_Xml0.Xnand0.MPMOS0_g N_VDD!_Xml0.Xnand0.MPMOS0_s
+ N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14
+ PD=1.37e-06 PS=1.26e-06
mXsl0.Xnor0.MPMOS1 XSL0.XNOR0.NET1 N_XSL0.N2_Xsl0.Xnor0.MPMOS1_g
+ N_VDD!_Xsl0.Xnor0.MPMOS1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=3.55e-07
+ AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXsl0.Xnor0.MPMOS0 N_XSL0.N3_Xsl0.Xnor0.MPMOS0_d N_RST_Xsl0.Xnor0.MPMOS0_g
+ XSL0.XNOR0.NET1 N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=3.55e-07
+ AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXml0.Xi0.MM0 N_XML0.N1_Xml0.Xi0.MM0_d N_D_Xml0.Xi0.MM0_g N_VSS!_Xml0.Xi0.MM0_s
+ N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14
+ PD=8.6e-07 PS=8.6e-07
mXml0.Xi0.MM1 N_XML0.N1_Xml0.Xi0.MM1_d N_D_Xml0.Xi0.MM1_g N_VDD!_Xml0.Xi0.MM1_s
+ N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14 AS=4.305e-14
+ PD=1.03e-06 PS=1.03e-06
mXml0.Xi1.MM0 N_N_Xml0.Xi1.MM0_d N_XML0.N2_Xml0.Xi1.MM0_g N_VSS!_Xml0.Xi1.MM0_s
+ N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14
+ PD=8.6e-07 PS=8.6e-07
mXml0.Xi1.MM1 N_N_Xml0.Xi1.MM1_d N_XML0.N2_Xml0.Xi1.MM1_g N_VDD!_Xml0.Xi1.MM1_s
+ N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14 AS=4.305e-14
+ PD=1.03e-06 PS=1.03e-06
mXsl0.Xi0.MM0 N_XSL0.N2_Xsl0.Xi0.MM0_d N_XSL0.N1_Xsl0.Xi0.MM0_g
+ N_VSS!_Xsl0.Xi0.MM0_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.25e-07
+ AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xi0.MM1 N_XSL0.N2_Xsl0.Xi0.MM1_d N_XSL0.N1_Xsl0.Xi0.MM1_g
+ N_VDD!_Xsl0.Xi0.MM1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=4.1e-07
+ AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXsl0.Xi1.MM0 N_Q_Xsl0.Xi1.MM0_d N_XSL0.N2_Xsl0.Xi1.MM0_g N_VSS!_Xsl0.Xi1.MM0_s
+ N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14
+ PD=8.6e-07 PS=8.6e-07
mXsl0.Xi1.MM1 N_Q_Xsl0.Xi1.MM1_d N_XSL0.N2_Xsl0.Xi1.MM1_g N_VDD!_Xsl0.Xi1.MM1_s
+ N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14 AS=4.305e-14
+ PD=1.03e-06 PS=1.03e-06
mXI0.MM0 N_CLKI_BAR_XI0.MM0_d N_CLK_XI0.MM0_g N_VSS!_XI0.MM0_s
+ N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14
+ PD=9e-07 PS=9e-07
mXI0.MM1 N_CLKI_BAR_XI0.MM1_d N_CLK_XI0.MM1_g N_VDD!_XI0.MM1_s N_VDD!_XI0.MM1_b
+ PMOS_VTG L=6e-08 W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06
+ PS=1.08e-06
mXI1.MM0 N_CLKI_XI1.MM0_d N_CLKI_BAR_XI1.MM0_g N_VSS!_XI1.MM0_s
+ N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14
+ PD=9e-07 PS=9e-07
mXI1.MM1 N_CLKI_XI1.MM1_d N_CLKI_BAR_XI1.MM1_g N_VDD!_XI1.MM1_s N_VDD!_XI0.MM1_b
+ PMOS_VTG L=6e-08 W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06
+ PS=1.08e-06
mXI2.MM0 N_RST_BAR_XI2.MM0_d N_RST_XI2.MM0_g N_VSS!_XI2.MM0_s
+ N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14
+ PD=9e-07 PS=9e-07
mXI2.MM1 N_RST_BAR_XI2.MM1_d N_RST_XI2.MM1_g N_VDD!_XI2.MM1_s N_VDD!_XI2.MM1_b
+ PMOS_VTG L=6e-08 W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06
+ PS=1.08e-06
mXml0.Xtg0.MM0 N_XML0.N1_Xml0.Xtg0.MM0_d N_CLKI_BAR_Xml0.Xtg0.MM0_g
+ N_XML0.N2_Xml0.Xtg0.MM0_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=2.65e-07
+ AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXml0.Xtg0.MM1 N_XML0.N1_Xml0.Xtg0.MM1_d N_CLKI_Xml0.Xtg0.MM1_g
+ N_XML0.N2_Xml0.Xtg0.MM1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=2.5e-07
+ AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXml0.Xtg1.MM0 N_XML0.N4_Xml0.Xtg1.MM0_d N_CLKI_Xml0.Xtg1.MM0_g
+ N_XML0.N2_Xml0.Xtg1.MM0_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=2.65e-07
+ AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXml0.Xtg1.MM1 N_XML0.N4_Xml0.Xtg1.MM1_d N_CLKI_BAR_Xml0.Xtg1.MM1_g
+ N_XML0.N2_Xml0.Xtg1.MM1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=2.5e-07
+ AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xtg1.MM0 N_N_Xsl0.Xtg1.MM0_d N_CLKI_Xsl0.Xtg1.MM0_g
+ N_XSL0.N1_Xsl0.Xtg1.MM0_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=2.65e-07
+ AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXsl0.Xtg1.MM1 N_N_Xsl0.Xtg1.MM1_d N_CLKI_BAR_Xsl0.Xtg1.MM1_g
+ N_XSL0.N1_Xsl0.Xtg1.MM1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=2.5e-07
+ AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xtg0.MM0 N_XSL0.N3_Xsl0.Xtg0.MM0_d N_CLKI_BAR_Xsl0.Xtg0.MM0_g
+ N_XSL0.N1_Xsl0.Xtg0.MM0_s N_VSS!_Xml0.Xi0.MM0_b NMOS_VTG L=6e-08 W=2.65e-07
+ AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXsl0.Xtg0.MM1 N_XSL0.N3_Xsl0.Xtg0.MM1_d N_CLKI_Xsl0.Xtg0.MM1_g
+ N_XSL0.N1_Xsl0.Xtg0.MM1_s N_VDD!_Xml0.Xi0.MM1_b PMOS_VTG L=6e-08 W=2.5e-07
+ AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
*
.include "DFSR.pex.netlist.DFSR.pxi"
*
.ends
*
*
.subckt loaded_flip_flop d rst q clk 
xdfsr0 clk d q rst DFSR
c0 q vss! 6e-15
.ends loaded_flip_flop
