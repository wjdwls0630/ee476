** Generated for: hspiceD
** Generated on: Nov 28 17:40:42 2021
** Design library name: cad6
** Design cell name: ALU_NAND_CELL_XOR
** Design view name: schematic
.GLOBAL vss! vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad6
** Cell name: MUX2_X1
** View name: schematic
.subckt MUX2_X1 a b s z
m_i_4 net_1 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_5 z_neg x1 net_1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_2 z_neg s net_0 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_3 net_0 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_10 vss! s x1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_6 net_2 s z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_8 vdd! a net_2 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_9 net_3 x1 z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_7 vdd! b net_3 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_11 vdd! s x1 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends MUX2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INV_X1
** View name: schematic
.subckt INV_X1 a zn
m_i_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INVMUX2_X1
** View name: schematic
.subckt INVMUX2_X1 a b s zn
xi0 a b s z MUX2_X1
xi1 z zn INV_X1
.ends INVMUX2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INVMUX4_X1
** View name: schematic
.subckt INVMUX4_X1 a b c d s<1> s<0> zn
xi2 net1 net2 s<1> zn INVMUX2_X1
xi1 c d s<0> net2 MUX2_X1
xi0 a b s<0> net1 MUX2_X1
.ends INVMUX4_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: NAND2_X1
** View name: schematic
.subckt NAND2_X1 a1 a2 zn
m_i_3 zn a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_2 vdd! a1 zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 zn a1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 net_0 a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends NAND2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: XNOR2_X1
** View name: schematic
.subckt XNOR2_X1 a b zn
m_i_48 net_003 a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_53 vdd! b net_003 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_29 net_000 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_36 vdd! b net_000 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_42 zn net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_0 net_001 a net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_5 vss! b net_001 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_11 net_002 net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_17 zn a net_002 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_23 net_002 b zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends XNOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: NOR2_X1
** View name: schematic
.subckt NOR2_X1 a1 a2 zn
m_i_1 zn a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 vss! a1 zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_2 zn a1 net_0 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_3 net_0 a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends NOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: LOGIC_UNIT
** View name: schematic
.subckt LOGIC_UNIT a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> b<15> b<14> b<13> b<12> b<11> b<10> b<9> b<8> b<7> b<6> b<5> b<4> b<3> b<2> b<1> b<0> logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> s<1> s<0>
xi0<15> nand<15> xnor<15> nor<15> a<15> s<1> s<0> logic_out<15> INVMUX4_X1
xi0<14> nand<14> xnor<14> nor<14> a<14> s<1> s<0> logic_out<14> INVMUX4_X1
xi0<13> nand<13> xnor<13> nor<13> a<13> s<1> s<0> logic_out<13> INVMUX4_X1
xi0<12> nand<12> xnor<12> nor<12> a<12> s<1> s<0> logic_out<12> INVMUX4_X1
xi0<11> nand<11> xnor<11> nor<11> a<11> s<1> s<0> logic_out<11> INVMUX4_X1
xi0<10> nand<10> xnor<10> nor<10> a<10> s<1> s<0> logic_out<10> INVMUX4_X1
xi0<9> nand<9> xnor<9> nor<9> a<9> s<1> s<0> logic_out<9> INVMUX4_X1
xi0<8> nand<8> xnor<8> nor<8> a<8> s<1> s<0> logic_out<8> INVMUX4_X1
xi0<7> nand<7> xnor<7> nor<7> a<7> s<1> s<0> logic_out<7> INVMUX4_X1
xi0<6> nand<6> xnor<6> nor<6> a<6> s<1> s<0> logic_out<6> INVMUX4_X1
xi0<5> nand<5> xnor<5> nor<5> a<5> s<1> s<0> logic_out<5> INVMUX4_X1
xi0<4> nand<4> xnor<4> nor<4> a<4> s<1> s<0> logic_out<4> INVMUX4_X1
xi0<3> nand<3> xnor<3> nor<3> a<3> s<1> s<0> logic_out<3> INVMUX4_X1
xi0<2> nand<2> xnor<2> nor<2> a<2> s<1> s<0> logic_out<2> INVMUX4_X1
xi0<1> nand<1> xnor<1> nor<1> a<1> s<1> s<0> logic_out<1> INVMUX4_X1
xi0<0> nand<0> xnor<0> nor<0> a<0> s<1> s<0> logic_out<0> INVMUX4_X1
xi1<15> a<15> b<15> nand<15> NAND2_X1
xi1<14> a<14> b<14> nand<14> NAND2_X1
xi1<13> a<13> b<13> nand<13> NAND2_X1
xi1<12> a<12> b<12> nand<12> NAND2_X1
xi1<11> a<11> b<11> nand<11> NAND2_X1
xi1<10> a<10> b<10> nand<10> NAND2_X1
xi1<9> a<9> b<9> nand<9> NAND2_X1
xi1<8> a<8> b<8> nand<8> NAND2_X1
xi1<7> a<7> b<7> nand<7> NAND2_X1
xi1<6> a<6> b<6> nand<6> NAND2_X1
xi1<5> a<5> b<5> nand<5> NAND2_X1
xi1<4> a<4> b<4> nand<4> NAND2_X1
xi1<3> a<3> b<3> nand<3> NAND2_X1
xi1<2> a<2> b<2> nand<2> NAND2_X1
xi1<1> a<1> b<1> nand<1> NAND2_X1
xi1<0> a<0> b<0> nand<0> NAND2_X1
xi2<15> a<15> b<15> xnor<15> XNOR2_X1
xi2<14> a<14> b<14> xnor<14> XNOR2_X1
xi2<13> a<13> b<13> xnor<13> XNOR2_X1
xi2<12> a<12> b<12> xnor<12> XNOR2_X1
xi2<11> a<11> b<11> xnor<11> XNOR2_X1
xi2<10> a<10> b<10> xnor<10> XNOR2_X1
xi2<9> a<9> b<9> xnor<9> XNOR2_X1
xi2<8> a<8> b<8> xnor<8> XNOR2_X1
xi2<7> a<7> b<7> xnor<7> XNOR2_X1
xi2<6> a<6> b<6> xnor<6> XNOR2_X1
xi2<5> a<5> b<5> xnor<5> XNOR2_X1
xi2<4> a<4> b<4> xnor<4> XNOR2_X1
xi2<3> a<3> b<3> xnor<3> XNOR2_X1
xi2<2> a<2> b<2> xnor<2> XNOR2_X1
xi2<1> a<1> b<1> xnor<1> XNOR2_X1
xi2<0> a<0> b<0> xnor<0> XNOR2_X1
xi3<15> a<15> b<15> nor<15> NOR2_X1
xi3<14> a<14> b<14> nor<14> NOR2_X1
xi3<13> a<13> b<13> nor<13> NOR2_X1
xi3<12> a<12> b<12> nor<12> NOR2_X1
xi3<11> a<11> b<11> nor<11> NOR2_X1
xi3<10> a<10> b<10> nor<10> NOR2_X1
xi3<9> a<9> b<9> nor<9> NOR2_X1
xi3<8> a<8> b<8> nor<8> NOR2_X1
xi3<7> a<7> b<7> nor<7> NOR2_X1
xi3<6> a<6> b<6> nor<6> NOR2_X1
xi3<5> a<5> b<5> nor<5> NOR2_X1
xi3<4> a<4> b<4> nor<4> NOR2_X1
xi3<3> a<3> b<3> nor<3> NOR2_X1
xi3<2> a<2> b<2> nor<2> NOR2_X1
xi3<1> a<1> b<1> nor<1> NOR2_X1
xi3<0> a<0> b<0> nor<0> NOR2_X1
.ends LOGIC_UNIT
** End of subcircuit definition.

** Library name: cad6
** Cell name: INV_X4
** View name: schematic
.subckt INV_X4 a zn
m_i_1_0_x4_0 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_1 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_2 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_3 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0_0_x4_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_1 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_2 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_3 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV_X4
** End of subcircuit definition.

** Library name: cad6
** Cell name: NOR4_X1
** View name: schematic
.subckt NOR4_X1 a1 a2 a3 a4 zn
m_i_2 vss! a3 zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_3 zn a4 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0 vss! a1 zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 zn a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_6 net_1 a3 net_2 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_7 net_2 a4 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_4 zn a1 net_0 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_5 net_0 a2 net_1 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
.ends NOR4_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: NAND4_X1
** View name: schematic
.subckt NAND4_X1 a1 a2 a3 a4 zn
m_i_6 vdd! a3 zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_7 zn a4 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_4 vdd! a1 zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_5 zn a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_2 net_1 a3 net_2 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_3 net_2 a4 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 zn a1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_1 net_0 a2 net_1 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
.ends NAND4_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: NAND3_X1
** View name: schematic
.subckt NAND3_X1 a1 a2 a3 zn
m_i_5 zn a3 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_3 zn a1 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_4 vdd! a2 zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_2 net_1 a3 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 zn a1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_1 net_0 a2 net_1 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
.ends NAND3_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: FA_X1
** View name: schematic
.subckt FA_X1 a b ci co s
m_instance_284 net_010 ci net_005 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_280 net_009 b net_010 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_275 vdd! a net_009 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_251 net_007 a net_001 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_246 vdd! b net_007 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_239 co net_001 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_instance_315 s net_005 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_269 net_008 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_263 vdd! b net_008 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_257 net_001 ci net_008 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_309 net_011 b vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_297 vdd! ci net_011 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_303 net_011 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_290 net_005 net_001 net_011 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_203 net_004 ci net_005 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_199 net_003 b net_004 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_194 vss! a net_003 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_159 co net_001 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_233 s net_005 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_166 vss! b net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_170 net_000 a net_001 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_176 net_001 ci net_002 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_209 net_005 net_001 net_006 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_215 vss! ci net_006 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_188 net_002 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_182 vss! b net_002 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_227 net_006 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_221 net_006 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
.ends FA_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: 4B_RCA
** View name: schematic
.subckt cad6_4B_RCA_schematic a<3> a<2> a<1> a<0> b<3> b<2> b<1> b<0> ci co s<3> s<2> s<1> s<0>
xi3 a<3> b<3> ci_3 co s<3> FA_X1
xi2 a<2> b<2> ci_2 ci_3 s<2> FA_X1
xi1 a<1> b<1> ci_1 ci_2 s<1> FA_X1
xi0 a<0> b<0> ci ci_1 s<0> FA_X1
.ends cad6_4B_RCA_schematic
** End of subcircuit definition.

** Library name: cad6
** Cell name: 4B_CSA
** View name: schematic
.subckt cad6_4B_CSA_schematic a<3> a<2> a<1> a<0> b<3> b<2> b<1> b<0> ci co s<3> s<2> s<1> s<0>
xi1 a<3> a<2> a<1> a<0> b<3> b<2> b<1> b<0> vdd! c_1 s_1<3> s_1<2> s_1<1> s_1<0> cad6_4B_RCA_schematic
xi0 a<3> a<2> a<1> a<0> b<3> b<2> b<1> b<0> vss! c_0 s_0<3> s_0<2> s_0<1> s_0<0> cad6_4B_RCA_schematic
xi3<3> s_0<3> s_1<3> ci s<3> MUX2_X1
xi3<2> s_0<2> s_1<2> ci s<2> MUX2_X1
xi3<1> s_0<1> s_1<1> ci s<1> MUX2_X1
xi3<0> s_0<0> s_1<0> ci s<0> MUX2_X1
xi2 c_0 c_1 ci co MUX2_X1
.ends cad6_4B_CSA_schematic
** End of subcircuit definition.

** Library name: cad6
** Cell name: 16B_CSA
** View name: schematic
.subckt cad6_16B_CSA_schematic a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> b<15> b<14> b<13> b<12> b<11> b<10> b<9> b<8> b<7> b<6> b<5> b<4> b<3> b<2> b<1> b<0> ci co s<15> s<14> s<13> s<12> s<11> s<10> s<9> s<8> s<7> s<6> s<5> s<4> s<3> s<2> s<1> s<0>
xi2 a<15> a<14> a<13> a<12> b<15> b<14> b<13> b<12> c_2 co s<15> s<14> s<13> s<12> cad6_4B_CSA_schematic
xi1 a<11> a<10> a<9> a<8> b<11> b<10> b<9> b<8> c_1 c_2 s<11> s<10> s<9> s<8> cad6_4B_CSA_schematic
xi0 a<7> a<6> a<5> a<4> b<7> b<6> b<5> b<4> c_0 c_1 s<7> s<6> s<5> s<4> cad6_4B_CSA_schematic
xi3 a<3> a<2> a<1> a<0> b<3> b<2> b<1> b<0> ci c_0 s<3> s<2> s<1> s<0> cad6_4B_RCA_schematic
.ends cad6_16B_CSA_schematic
** End of subcircuit definition.

** Library name: cad6
** Cell name: NAND_CELL_XOR2_X1
** View name: schematic
.subckt NAND_CELL_XOR2_X1 a b z
m_i_30 net_002 a net_000 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_35 vdd! b net_002 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_41 net_003 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_47 z a net_003 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_53 net_003 b z vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_19 net_001 a z vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_24 vss! b net_001 vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 net_000 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_13 z net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_7 vss! b net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends NAND_CELL_XOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: ARITMETIC_UNIT_NAND_XOR
** View name: schematic
.subckt ARITMETIC_UNIT_NAND_XOR a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> aritmetic_out<15> aritmetic_out<14> aritmetic_out<13> aritmetic_out<12> aritmetic_out<11> aritmetic_out<10> aritmetic_out<9> aritmetic_out<8> aritmetic_out<7> aritmetic_out<6> aritmetic_out<5> aritmetic_out<4> aritmetic_out<3> aritmetic_out<2> aritmetic_out<1> aritmetic_out<0> a_temp<15> b<15> b<14> b<13> b<12> b<11> b<10> b<9> b<8> b<7> b<6> b<5> b<4> b<3> b<2> b<1> b<0> co s
xi0 a_temp<15> a_temp<14> a_temp<13> a_temp<12> a_temp<11> a_temp<10> a_temp<9> a_temp<8> a_temp<7> a_temp<6> a_temp<5> a_temp<4> a_temp<3> a_temp<2> a_temp<1> a_temp<0> b<15> b<14> b<13> b<12> b<11> b<10> b<9> b<8> b<7> b<6> b<5> b<4> b<3> b<2> b<1> b<0> s co aritmetic_out<15> aritmetic_out<14> aritmetic_out<13> aritmetic_out<12> aritmetic_out<11> aritmetic_out<10> aritmetic_out<9> aritmetic_out<8> aritmetic_out<7> aritmetic_out<6> aritmetic_out<5> aritmetic_out<4> aritmetic_out<3> aritmetic_out<2> aritmetic_out<1> aritmetic_out<0> cad6_16B_CSA_schematic
xi3<15> a<15> s a_temp<15> NAND_CELL_XOR2_X1
xi3<14> a<14> s a_temp<14> NAND_CELL_XOR2_X1
xi3<13> a<13> s a_temp<13> NAND_CELL_XOR2_X1
xi3<12> a<12> s a_temp<12> NAND_CELL_XOR2_X1
xi3<11> a<11> s a_temp<11> NAND_CELL_XOR2_X1
xi3<10> a<10> s a_temp<10> NAND_CELL_XOR2_X1
xi3<9> a<9> s a_temp<9> NAND_CELL_XOR2_X1
xi3<8> a<8> s a_temp<8> NAND_CELL_XOR2_X1
xi3<7> a<7> s a_temp<7> NAND_CELL_XOR2_X1
xi3<6> a<6> s a_temp<6> NAND_CELL_XOR2_X1
xi3<5> a<5> s a_temp<5> NAND_CELL_XOR2_X1
xi3<4> a<4> s a_temp<4> NAND_CELL_XOR2_X1
xi3<3> a<3> s a_temp<3> NAND_CELL_XOR2_X1
xi3<2> a<2> s a_temp<2> NAND_CELL_XOR2_X1
xi3<1> a<1> s a_temp<1> NAND_CELL_XOR2_X1
xi3<0> a<0> s a_temp<0> NAND_CELL_XOR2_X1
.ends ARITMETIC_UNIT_NAND_XOR
** End of subcircuit definition.

** Library name: cad6
** Cell name: ALU_NAND_CELL_XOR
** View name: schematic
xi0 op0<15> op0<14> op0<13> op0<12> op0<11> op0<10> op0<9> op0<8> op0<7> op0<6> op0<5> op0<4> op0<3> op0<2> op0<1> op0<0> op1<15> op1<14> op1<13> op1<12> op1<11> op1<10> op1<9> op1<8> op1<7> op1<6> op1<5> op1<4> op1<3> op1<2> op1<1> op1<0> logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> ctrl<1> ctrl<0> LOGIC_UNIT
xi3<15> logic_out<15> aritmetic_out<15> ctrl<2> alu_pre<15> MUX2_X1
xi3<14> logic_out<14> aritmetic_out<14> ctrl<2> alu_pre<14> MUX2_X1
xi3<13> logic_out<13> aritmetic_out<13> ctrl<2> alu_pre<13> MUX2_X1
xi3<12> logic_out<12> aritmetic_out<12> ctrl<2> alu_pre<12> MUX2_X1
xi3<11> logic_out<11> aritmetic_out<11> ctrl<2> alu_pre<11> MUX2_X1
xi3<10> logic_out<10> aritmetic_out<10> ctrl<2> alu_pre<10> MUX2_X1
xi3<9> logic_out<9> aritmetic_out<9> ctrl<2> alu_pre<9> MUX2_X1
xi3<8> logic_out<8> aritmetic_out<8> ctrl<2> alu_pre<8> MUX2_X1
xi3<7> logic_out<7> aritmetic_out<7> ctrl<2> alu_pre<7> MUX2_X1
xi3<6> logic_out<6> aritmetic_out<6> ctrl<2> alu_pre<6> MUX2_X1
xi3<5> logic_out<5> aritmetic_out<5> ctrl<2> alu_pre<5> MUX2_X1
xi3<4> logic_out<4> aritmetic_out<4> ctrl<2> alu_pre<4> MUX2_X1
xi3<3> logic_out<3> aritmetic_out<3> ctrl<2> alu_pre<3> MUX2_X1
xi3<2> logic_out<2> aritmetic_out<2> ctrl<2> alu_pre<2> MUX2_X1
xi3<1> logic_out<1> aritmetic_out<1> ctrl<2> alu_pre<1> MUX2_X1
xi3<0> logic_out<0> aritmetic_out<0> ctrl<2> alu_pre<0> MUX2_X1
xi7 c0n c_flag INV_X4
xi21 zflag_inv z_flag INV_X4
xi9 pf n_flag INV_X4
xi4<15> alu_inv<15> alu_out<15> INV_X4
xi4<14> alu_inv<14> alu_out<14> INV_X4
xi4<13> alu_inv<13> alu_out<13> INV_X4
xi4<12> alu_inv<12> alu_out<12> INV_X4
xi4<11> alu_inv<11> alu_out<11> INV_X4
xi4<10> alu_inv<10> alu_out<10> INV_X4
xi4<9> alu_inv<9> alu_out<9> INV_X4
xi4<8> alu_inv<8> alu_out<8> INV_X4
xi4<7> alu_inv<7> alu_out<7> INV_X4
xi4<6> alu_inv<6> alu_out<6> INV_X4
xi4<5> alu_inv<5> alu_out<5> INV_X4
xi4<4> alu_inv<4> alu_out<4> INV_X4
xi4<3> alu_inv<3> alu_out<3> INV_X4
xi4<2> alu_inv<2> alu_out<2> INV_X4
xi4<1> alu_inv<1> alu_out<1> INV_X4
xi4<0> alu_inv<0> alu_out<0> INV_X4
xi6 co c0n INV_X1
xi20 aritmetic_out<15> aritmetic_out_15_n INV_X1
xi19 op1<15> op1_15_n INV_X1
xi18 a_temp a_temp_n INV_X1
xi8 alu_pre<15> pf INV_X1
xi5<15> alu_pre<15> alu_inv<15> INV_X1
xi5<14> alu_pre<14> alu_inv<14> INV_X1
xi5<13> alu_pre<13> alu_inv<13> INV_X1
xi5<12> alu_pre<12> alu_inv<12> INV_X1
xi5<11> alu_pre<11> alu_inv<11> INV_X1
xi5<10> alu_pre<10> alu_inv<10> INV_X1
xi5<9> alu_pre<9> alu_inv<9> INV_X1
xi5<8> alu_pre<8> alu_inv<8> INV_X1
xi5<7> alu_pre<7> alu_inv<7> INV_X1
xi5<6> alu_pre<6> alu_inv<6> INV_X1
xi5<5> alu_pre<5> alu_inv<5> INV_X1
xi5<4> alu_pre<4> alu_inv<4> INV_X1
xi5<3> alu_pre<3> alu_inv<3> INV_X1
xi5<2> alu_pre<2> alu_inv<2> INV_X1
xi5<1> alu_pre<1> alu_inv<1> INV_X1
xi5<0> alu_pre<0> alu_inv<0> INV_X1
xi13 alu_pre<3> alu_pre<2> alu_pre<1> alu_pre<0> z3 NOR4_X1
xi12 alu_pre<7> alu_pre<6> alu_pre<5> alu_pre<4> z2 NOR4_X1
xi11 alu_pre<11> alu_pre<10> alu_pre<9> alu_pre<8> z1 NOR4_X1
xi10 alu_pre<15> alu_pre<14> alu_pre<13> alu_pre<12> z0 NOR4_X1
xi14 z0 z1 z2 z3 zflag_inv NAND4_X1
xi16 a_temp_n op1_15_n aritmetic_out<15> ov1 NAND3_X1
xi15 a_temp op1<15> aritmetic_out_15_n ov0 NAND3_X1
xi17 ov0 ov1 v_flag NAND2_X1
xi1 op0<15> op0<14> op0<13> op0<12> op0<11> op0<10> op0<9> op0<8> op0<7> op0<6> op0<5> op0<4> op0<3> op0<2> op0<1> op0<0> aritmetic_out<15> aritmetic_out<14> aritmetic_out<13> aritmetic_out<12> aritmetic_out<11> aritmetic_out<10> aritmetic_out<9> aritmetic_out<8> aritmetic_out<7> aritmetic_out<6> aritmetic_out<5> aritmetic_out<4> aritmetic_out<3> aritmetic_out<2> aritmetic_out<1> aritmetic_out<0> a_temp op1<15> op1<14> op1<13> op1<12> op1<11> op1<10> op1<9> op1<8> op1<7> op1<6> op1<5> op1<4> op1<3> op1<2> op1<1> op1<0> co ctrl<0> ARITMETIC_UNIT_NAND_XOR
.END
