.GLOBAL vdd! vss!


.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2

* File: DFSR.pex.netlist
* Created: Sun Nov  7 21:57:51 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.subckt DFSR CLK D Q RST 
* 
mXml0.Xnand0.MNMOS1 XML0.XNAND0.NET2 N VSS! VSS! NMOS_VTG L=6e-08 W=2.5e-07
+ AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXml0.Xnand0.MNMOS0 XML0.N4 RST_BAR XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08
+ W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXsl0.Xnor0.MNMOS1 XSL0.N3 XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08 W=9.5e-08
+ AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXsl0.Xnor0.MNMOS0 XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08 W=9.5e-08 AD=1.52e-14
+ AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXml0.Xnand0.MPMOS1 XML0.N4 N VDD! VDD! PMOS_VTG L=6e-08 W=5.25e-07 AD=8.4e-14
+ AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXml0.Xnand0.MPMOS0 XML0.N4 RST_BAR VDD! VDD! PMOS_VTG L=6e-08 W=5.25e-07
+ AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXsl0.Xnor0.MPMOS1 XSL0.XNOR0.NET1 XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08 W=3.55e-07
+ AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXsl0.Xnor0.MPMOS0 XSL0.N3 RST XSL0.XNOR0.NET1 VDD! PMOS_VTG L=6e-08 W=3.55e-07
+ AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXI0.MM0 CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07 AD=3.6225e-14
+ AS=3.6225e-14 PD=9e-07 PS=9e-07
mXI0.MM1 CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07 AD=4.5675e-14
+ AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXI1.MM0 CLKI CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07 AD=3.6225e-14
+ AS=3.6225e-14 PD=9e-07 PS=9e-07
mXI1.MM1 CLKI CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07 AD=4.5675e-14
+ AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXI2.MM0 RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07 AD=3.6225e-14
+ AS=3.6225e-14 PD=9e-07 PS=9e-07
mXI2.MM1 RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07 AD=4.5675e-14
+ AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXml0.Xi0.MM0 XML0.N1 D VSS! VSS! NMOS_VTG L=6e-08 W=3.25e-07 AD=3.4125e-14
+ AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXml0.Xi0.MM1 XML0.N1 D VDD! VDD! PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14
+ AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXml0.Xi1.MM0 N XML0.N2 VSS! VSS! NMOS_VTG L=6e-08 W=3.25e-07 AD=3.4125e-14
+ AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXml0.Xi1.MM1 N XML0.N2 VDD! VDD! PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14
+ AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXsl0.Xi0.MM0 XSL0.N2 XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08 W=3.25e-07
+ AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xi0.MM1 XSL0.N2 XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14
+ AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXsl0.Xi1.MM0 Q XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08 W=3.25e-07 AD=3.4125e-14
+ AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xi1.MM1 Q XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08 W=4.1e-07 AD=4.305e-14
+ AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXml0.Xtg0.MM0 XML0.N1 CLKI_BAR XML0.N2 VSS! NMOS_VTG L=6e-08 W=2.65e-07
+ AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXml0.Xtg0.MM1 XML0.N1 CLKI XML0.N2 VDD! PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14
+ AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXml0.Xtg1.MM0 XML0.N4 CLKI XML0.N2 VSS! NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14
+ AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXml0.Xtg1.MM1 XML0.N4 CLKI_BAR XML0.N2 VDD! PMOS_VTG L=6e-08 W=2.5e-07
+ AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xtg1.MM0 N CLKI XSL0.N1 VSS! NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14
+ AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXsl0.Xtg1.MM1 N CLKI_BAR XSL0.N1 VDD! PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14
+ AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXsl0.Xtg0.MM0 XSL0.N3 CLKI_BAR XSL0.N1 VSS! NMOS_VTG L=6e-08 W=2.65e-07
+ AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXsl0.Xtg0.MM1 XSL0.N3 CLKI XSL0.N1 VDD! PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14
+ AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
c_9 N 0 0.159231f
c_21 RST_BAR 0 0.189728f
c_28 RST 0 0.191671f
c_42 CLKI_BAR 0 0.368607f
c_49 XML0.N1 0 0.0382055f
c_57 XML0.N2 0 0.127547f
c_65 XML0.N4 0 0.0452973f
c_74 XSL0.N1 0 0.12236f
c_84 XSL0.N2 0 0.194773f
c_94 XSL0.N3 0 0.0533432f
c_110 VSS! 0 0.408952f
c_126 VDD! 0 0.43723f
c_139 CLKI 0 0.29199f
c_143 CLK 0 0.100368f
c_149 D 0 0.0873897f
c_156 Q 0 0.0180042f
*
.include "DFSR.pex.netlist.DFSR.pxi"
*
.ends
*
*

.subckt loaded_flip_flop d rst q clk 
xdfsr0 clk d q rst DFSR
c0 q vss! 6e-15
.ends loaded_flip_flop
