

.OPTION

.subckt rc_series vi vo
r0 vi vo 1e3
c1 vo 0 1e-12
.ends rc_series
.END
