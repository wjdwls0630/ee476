* File: /mmfs1/home/jarenas/ee476/jarenas_git/cad6/netlist/PEX/ALU.pex.netlist
* Created: Wed Dec  8 23:52:41 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.GLOBAL vss! vdd!


.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2

.subckt ALU
+ alu_out<0> alu_out<1> alu_out<2> alu_out<3> alu_out<4> alu_out<5> alu_out<6> alu_out<7>
+ alu_out<8> alu_out<9> alu_out<10> alu_out<11> alu_out<12> alu_out<13> alu_out<14> alu_out<15>
+ op0<0> op0<1> op0<2> op0<3> op0<4> op0<5> op0<6> op0<7>
+ op0<8> op0<9> op0<10> op0<11> op0<12> op0<13> op0<14> op0<15>
+ op1<0> op1<1> op1<2> op1<3> op1<4> op1<5> op1<6> op1<7>
+ op1<8> op1<9> op1<10> op1<11> op1<12> op1<13> op1<14> op1<15>
+ c_flag n_flag v_flag
+ ctrl<0> ctrl<1> ctrl<2>
* 
mXI17/MM_i_1__m0_m2__m0 VSS! OV1 XI17/NET_0__M0__M0 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI17/MM_i_0__m0_m2__m0 XI17/NET_0__M0__M0 OV0 V_FLAG VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI17/MM_i_0__m0_m2__m1 XI17/NET_0__M0__M1 OV0 V_FLAG VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI17/MM_i_1__m0_m2__m1 VSS! OV1 XI17/NET_0__M0__M1 VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI17/MM_i_3__m0_x2__m0 VDD! OV1 V_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI17/MM_i_2__m0_x2__m0 V_FLAG OV0 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI17/MM_i_2__m0_x2__m1 V_FLAG OV0 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI17/MM_i_3__m0_x2__m1 VDD! OV1 V_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI33/MM_i_0 CO_N CO VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI33/MM_i_1 CO_N CO VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI19/MM_i_0 OP1_N<15> OP1<15> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI19/MM_i_1 OP1_N<15> OP1<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI18/MM_i_0 OP0_TEMP_N<15> OP0_TEMP<15> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI18/MM_i_1 OP0_TEMP_N<15> OP0_TEMP<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI35/MM_i_0 ALU_PRE_N<15> ALU_PRE<15> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI35/MM_i_1 ALU_PRE_N<15> ALU_PRE<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI36/MM_i_0_0_x4_0 VSS! ALU_PRE_N<15> N_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI36/MM_i_0_0_x4_1 VSS! ALU_PRE_N<15> N_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI36/MM_i_0_0_x4_2 VSS! ALU_PRE_N<15> N_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI36/MM_i_0_0_x4_3 VSS! ALU_PRE_N<15> N_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI36/MM_i_1_0_x4_0 VDD! ALU_PRE_N<15> N_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI36/MM_i_1_0_x4_1 VDD! ALU_PRE_N<15> N_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI36/MM_i_1_0_x4_2 VDD! ALU_PRE_N<15> N_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI36/MM_i_1_0_x4_3 VDD! ALU_PRE_N<15> N_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI39<1>/MM_i_0 C0X<1> CTRL<1> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI39<1>/MM_i_1 C0X<1> CTRL<1> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI40<1>/MM_i_0_0_x4_0 VSS! C0X<1> CTRL_BUFF<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI40<1>/MM_i_0_0_x4_1 VSS! C0X<1> CTRL_BUFF<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI40<1>/MM_i_0_0_x4_2 VSS! C0X<1> CTRL_BUFF<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI40<1>/MM_i_0_0_x4_3 VSS! C0X<1> CTRL_BUFF<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI40<1>/MM_i_1_0_x4_0 VDD! C0X<1> CTRL_BUFF<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI40<1>/MM_i_1_0_x4_1 VDD! C0X<1> CTRL_BUFF<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI40<1>/MM_i_1_0_x4_2 VDD! C0X<1> CTRL_BUFF<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI40<1>/MM_i_1_0_x4_3 VDD! C0X<1> CTRL_BUFF<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI39<0>/MM_i_0 C0X<0> CTRL<0> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI39<0>/MM_i_1 C0X<0> CTRL<0> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI40<0>/MM_i_0_0_x4_0 VSS! C0X<0> CTRL_BUFF<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI40<0>/MM_i_0_0_x4_1 VSS! C0X<0> CTRL_BUFF<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI40<0>/MM_i_0_0_x4_2 VSS! C0X<0> CTRL_BUFF<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI40<0>/MM_i_0_0_x4_3 VSS! C0X<0> CTRL_BUFF<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI40<0>/MM_i_1_0_x4_0 VDD! C0X<0> CTRL_BUFF<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI40<0>/MM_i_1_0_x4_1 VDD! C0X<0> CTRL_BUFF<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI40<0>/MM_i_1_0_x4_2 VDD! C0X<0> CTRL_BUFF<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI40<0>/MM_i_1_0_x4_3 VDD! C0X<0> CTRL_BUFF<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI20/MM_i_0 ARITHMETIC_OUT_N<15> ARITHMETIC_OUT<15> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI20/MM_i_1 ARITHMETIC_OUT_N<15> ARITHMETIC_OUT<15> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI34/MM_i_0_0_x4_0 VSS! CO_N C_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI34/MM_i_0_0_x4_1 VSS! CO_N C_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI34/MM_i_0_0_x4_2 VSS! CO_N C_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI34/MM_i_0_0_x4_3 VSS! CO_N C_FLAG VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI34/MM_i_1_0_x4_0 VDD! CO_N C_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI34/MM_i_1_0_x4_1 VDD! CO_N C_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI34/MM_i_1_0_x4_2 VDD! CO_N C_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI34/MM_i_1_0_x4_3 VDD! CO_N C_FLAG VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI39<2>/MM_i_0 C0X<2> CTRL<2> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI39<2>/MM_i_1 C0X<2> CTRL<2> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI40<2>/MM_i_0_0_x4_0 VSS! C0X<2> CTRL_BUFF<2> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI40<2>/MM_i_0_0_x4_1 VSS! C0X<2> CTRL_BUFF<2> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI40<2>/MM_i_0_0_x4_2 VSS! C0X<2> CTRL_BUFF<2> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI40<2>/MM_i_0_0_x4_3 VSS! C0X<2> CTRL_BUFF<2> VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI40<2>/MM_i_1_0_x4_0 VDD! C0X<2> CTRL_BUFF<2> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI40<2>/MM_i_1_0_x4_1 VDD! C0X<2> CTRL_BUFF<2> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI40<2>/MM_i_1_0_x4_2 VDD! C0X<2> CTRL_BUFF<2> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI40<2>/MM_i_1_0_x4_3 VDD! C0X<2> CTRL_BUFF<2> VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI16/MM_i_2 XI16/NET_1 ARITHMETIC_OUT<15> VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI16/MM_i_1 XI16/NET_0 OP1_N<15> XI16/NET_1 VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI16/MM_i_0 OV1 OP0_TEMP_N<15> XI16/NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI16/MM_i_5 OV1 ARITHMETIC_OUT<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI16/MM_i_4 VDD! OP1_N<15> OV1 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI16/MM_i_3 OV1 OP0_TEMP_N<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI15/MM_i_2 XI15/NET_1 ARITHMETIC_OUT_N<15> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI15/MM_i_1 XI15/NET_0 OP1<15> XI15/NET_1 VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI15/MM_i_0 OV0 OP0_TEMP<15> XI15/NET_0 VSS! NMOS_VTL L=5e-08 W=4.15e-07
+ AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI15/MM_i_5 OV0 ARITHMETIC_OUT_N<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07
+ AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI15/MM_i_4 VDD! OP1<15> OV0 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI15/MM_i_3 OV0 OP0_TEMP<15> VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<15>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<0> ALU_OUT<15> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<15>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<0> ALU_OUT<15> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<15>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<0> ALU_OUT<15> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<15>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<0> ALU_OUT<15> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<15>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<0> ALU_OUT<15> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<15>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<0> ALU_OUT<15> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<15>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<0> ALU_OUT<15> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<15>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<0> ALU_OUT<15> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<15>/MM_i_0 XI31/XI2/NET3<0> ALU_PRE<15> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<15>/MM_i_1 XI31/XI2/NET3<0> ALU_PRE<15> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<15>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<15>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<15>/MM_i_4 XI31/XI2/XI0<15>/NET_1 XI31/LOGIC_OUT<15> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<15>/MM_i_5 XI31/XI2/XI0<15>/Z_NEG XI31/XI2/XI0<15>/X1
+ XI31/XI2/XI0<15>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<15>/MM_i_2 XI31/XI2/XI0<15>/Z_NEG CTRL_BUFF<2>
+ XI31/XI2/XI0<15>/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<15>/MM_i_3 XI31/XI2/XI0<15>/NET_0 ARITHMETIC_OUT<15> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<15>/MM_i_0 ALU_PRE<15> XI31/XI2/XI0<15>/Z_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<15>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<15>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<15>/MM_i_8 VDD! XI31/LOGIC_OUT<15> XI31/XI2/XI0<15>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<15>/MM_i_6 XI31/XI2/XI0<15>/NET_2 CTRL_BUFF<2>
+ XI31/XI2/XI0<15>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<15>/MM_i_9 XI31/XI2/XI0<15>/NET_3 XI31/XI2/XI0<15>/X1
+ XI31/XI2/XI0<15>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<15>/MM_i_7 VDD! ARITHMETIC_OUT<15> XI31/XI2/XI0<15>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<15>/MM_i_1 ALU_PRE<15> XI31/XI2/XI0<15>/Z_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI0/XI0/MM_i_1 XI31/XI0/XI0/XI0/NET_0 OP0<15> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI0/XI0/MM_i_0 XI31/XI0/XI0/NAND_OUT OP1<15> XI31/XI0/XI0/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI0/XI1/MM_i_0 XI31/XI0/XI0/XI1/NET_001 OP1<15>
+ XI31/XI0/XI0/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI0/XI1/MM_i_5 VSS! OP0<15> XI31/XI0/XI0/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI0/XI1/MM_i_11 XI31/XI0/XI0/XI1/NET_002 XI31/XI0/XI0/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI0/XI1/MM_i_17 XI31/XI0/XI0/XNOR_OUT OP1<15> XI31/XI0/XI0/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI0/XI1/MM_i_23 XI31/XI0/XI0/XI1/NET_002 OP0<15> XI31/XI0/XI0/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI0/XI2/MM_i_1 XI31/XI0/XI0/NOR_OUT OP0<15> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI0/XI2/MM_i_0 VSS! OP1<15> XI31/XI0/XI0/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI0/XI0/MM_i_3 XI31/XI0/XI0/NAND_OUT OP0<15> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI0/XI0/MM_i_2 VDD! OP1<15> XI31/XI0/XI0/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI0/XI1/MM_i_29 XI31/XI0/XI0/XI1/NET_000 OP1<15> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI0/XI1/MM_i_36 VDD! OP0<15> XI31/XI0/XI0/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI0/XI1/MM_i_42 XI31/XI0/XI0/XNOR_OUT XI31/XI0/XI0/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI0/XI1/MM_i_48 XI31/XI0/XI0/XI1/NET_003 OP1<15> XI31/XI0/XI0/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI0/XI1/MM_i_53 VDD! OP0<15> XI31/XI0/XI0/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI0/XI2/MM_i_3 XI31/XI0/XI0/XI2/NET_0 OP0<15> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI0/XI2/MM_i_2 XI31/XI0/XI0/NOR_OUT OP1<15> XI31/XI0/XI0/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI0/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<15> XI31/XI0/XI0/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI0/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<15> XI31/XI0/XI0/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI0/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI0/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI0/XI4/MM_i_4 XI31/XI0/XI0/XI4/NET_1 XI31/XI0/XI0/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI4/MM_i_5 XI31/XI0/XI0/XI4/Z_NEG XI31/XI0/XI0/XI4/X1
+ XI31/XI0/XI0/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI4/MM_i_2 XI31/XI0/XI0/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI0/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI4/MM_i_3 XI31/XI0/XI0/XI4/NET_0 OP0<15> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI0/XI4/MM_i_0 XI31/XI0/XI0/MUX1 XI31/XI0/XI0/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI0/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI0/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI0/XI4/MM_i_8 VDD! XI31/XI0/XI0/NOR_OUT XI31/XI0/XI0/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI4/MM_i_6 XI31/XI0/XI0/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI0/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI4/MM_i_9 XI31/XI0/XI0/XI4/NET_3 XI31/XI0/XI0/XI4/X1
+ XI31/XI0/XI0/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI4/MM_i_7 VDD! OP0<15> XI31/XI0/XI0/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI0/XI4/MM_i_1 XI31/XI0/XI0/MUX1 XI31/XI0/XI0/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI0/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI0/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_4 XI31/XI0/XI0/XI5/XI0/NET_1 XI31/XI0/XI0/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_5 XI31/XI0/XI0/XI5/XI0/Z_NEG XI31/XI0/XI0/XI5/XI0/X1
+ XI31/XI0/XI0/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_2 XI31/XI0/XI0/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI0/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_3 XI31/XI0/XI0/XI5/XI0/NET_0 XI31/XI0/XI0/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI0/XI5/XI0/MM_i_0 XI31/XI0/XI0/XI5/Z XI31/XI0/XI0/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI0/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI0/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI0/MUX0 XI31/XI0/XI0/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_6 XI31/XI0/XI0/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI0/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_9 XI31/XI0/XI0/XI5/XI0/NET_3 XI31/XI0/XI0/XI5/XI0/X1
+ XI31/XI0/XI0/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI0/MUX1 XI31/XI0/XI0/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI0/XI5/XI0/MM_i_1 XI31/XI0/XI0/XI5/Z XI31/XI0/XI0/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI0/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI0/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI0/XI3/MM_i_4 XI31/XI0/XI0/XI3/NET_1 XI31/XI0/XI0/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI3/MM_i_5 XI31/XI0/XI0/XI3/Z_NEG XI31/XI0/XI0/XI3/X1
+ XI31/XI0/XI0/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI3/MM_i_2 XI31/XI0/XI0/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI0/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI0/XI3/MM_i_3 XI31/XI0/XI0/XI3/NET_0 XI31/XI0/XI0/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI0/XI3/MM_i_0 XI31/XI0/XI0/MUX0 XI31/XI0/XI0/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI0/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI0/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI0/XI3/MM_i_8 VDD! XI31/XI0/XI0/NAND_OUT XI31/XI0/XI0/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI3/MM_i_6 XI31/XI0/XI0/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI0/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI3/MM_i_9 XI31/XI0/XI0/XI3/NET_3 XI31/XI0/XI0/XI3/X1
+ XI31/XI0/XI0/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI0/XI3/MM_i_7 VDD! XI31/XI0/XI0/XNOR_OUT XI31/XI0/XI0/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI0/XI3/MM_i_1 XI31/XI0/XI0/MUX0 XI31/XI0/XI0/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<14>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<1> ALU_OUT<14> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<14>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<1> ALU_OUT<14> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<14>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<1> ALU_OUT<14> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<14>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<1> ALU_OUT<14> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<14>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<1> ALU_OUT<14> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<14>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<1> ALU_OUT<14> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<14>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<1> ALU_OUT<14> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<14>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<1> ALU_OUT<14> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<14>/MM_i_0 XI31/XI2/NET3<1> XI31/XI2/ALU_PRE<14> VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI2/XI1<14>/MM_i_1 XI31/XI2/NET3<1> XI31/XI2/ALU_PRE<14> VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<14>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<14>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<14>/MM_i_4 XI31/XI2/XI0<14>/NET_1 XI31/LOGIC_OUT<14> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<14>/MM_i_5 XI31/XI2/XI0<14>/Z_NEG XI31/XI2/XI0<14>/X1
+ XI31/XI2/XI0<14>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<14>/MM_i_2 XI31/XI2/XI0<14>/Z_NEG CTRL_BUFF<2>
+ XI31/XI2/XI0<14>/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<14>/MM_i_3 XI31/XI2/XI0<14>/NET_0 XI31/ARITHMETIC_OUT<14> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<14>/MM_i_0 XI31/XI2/ALU_PRE<14> XI31/XI2/XI0<14>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<14>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<14>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<14>/MM_i_8 VDD! XI31/LOGIC_OUT<14> XI31/XI2/XI0<14>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<14>/MM_i_6 XI31/XI2/XI0<14>/NET_2 CTRL_BUFF<2>
+ XI31/XI2/XI0<14>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<14>/MM_i_9 XI31/XI2/XI0<14>/NET_3 XI31/XI2/XI0<14>/X1
+ XI31/XI2/XI0<14>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<14>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<14> XI31/XI2/XI0<14>/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI2/XI0<14>/MM_i_1 XI31/XI2/ALU_PRE<14> XI31/XI2/XI0<14>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI4/XI0/MM_i_1 XI31/XI0/XI4/XI0/NET_0 OP0<14> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI4/XI0/MM_i_0 XI31/XI0/XI4/NAND_OUT OP1<14> XI31/XI0/XI4/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI4/XI1/MM_i_0 XI31/XI0/XI4/XI1/NET_001 OP1<14>
+ XI31/XI0/XI4/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI4/XI1/MM_i_5 VSS! OP0<14> XI31/XI0/XI4/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI4/XI1/MM_i_11 XI31/XI0/XI4/XI1/NET_002 XI31/XI0/XI4/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI4/XI1/MM_i_17 XI31/XI0/XI4/XNOR_OUT OP1<14> XI31/XI0/XI4/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI4/XI1/MM_i_23 XI31/XI0/XI4/XI1/NET_002 OP0<14> XI31/XI0/XI4/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI4/XI2/MM_i_1 XI31/XI0/XI4/NOR_OUT OP0<14> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI4/XI2/MM_i_0 VSS! OP1<14> XI31/XI0/XI4/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI4/XI0/MM_i_3 XI31/XI0/XI4/NAND_OUT OP0<14> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI4/XI0/MM_i_2 VDD! OP1<14> XI31/XI0/XI4/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI4/XI1/MM_i_29 XI31/XI0/XI4/XI1/NET_000 OP1<14> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI4/XI1/MM_i_36 VDD! OP0<14> XI31/XI0/XI4/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI4/XI1/MM_i_42 XI31/XI0/XI4/XNOR_OUT XI31/XI0/XI4/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI4/XI1/MM_i_48 XI31/XI0/XI4/XI1/NET_003 OP1<14> XI31/XI0/XI4/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI4/XI1/MM_i_53 VDD! OP0<14> XI31/XI0/XI4/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI4/XI2/MM_i_3 XI31/XI0/XI4/XI2/NET_0 OP0<14> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI4/XI2/MM_i_2 XI31/XI0/XI4/NOR_OUT OP1<14> XI31/XI0/XI4/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI4/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<14> XI31/XI0/XI4/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI4/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<14> XI31/XI0/XI4/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI4/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI4/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI4/XI4/MM_i_4 XI31/XI0/XI4/XI4/NET_1 XI31/XI0/XI4/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI4/MM_i_5 XI31/XI0/XI4/XI4/Z_NEG XI31/XI0/XI4/XI4/X1
+ XI31/XI0/XI4/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI4/MM_i_2 XI31/XI0/XI4/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI4/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI4/MM_i_3 XI31/XI0/XI4/XI4/NET_0 OP0<14> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI4/XI4/MM_i_0 XI31/XI0/XI4/MUX1 XI31/XI0/XI4/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI4/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI4/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI4/XI4/MM_i_8 VDD! XI31/XI0/XI4/NOR_OUT XI31/XI0/XI4/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI4/MM_i_6 XI31/XI0/XI4/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI4/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI4/MM_i_9 XI31/XI0/XI4/XI4/NET_3 XI31/XI0/XI4/XI4/X1
+ XI31/XI0/XI4/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI4/MM_i_7 VDD! OP0<14> XI31/XI0/XI4/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI4/XI4/MM_i_1 XI31/XI0/XI4/MUX1 XI31/XI0/XI4/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI4/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI4/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_4 XI31/XI0/XI4/XI5/XI0/NET_1 XI31/XI0/XI4/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_5 XI31/XI0/XI4/XI5/XI0/Z_NEG XI31/XI0/XI4/XI5/XI0/X1
+ XI31/XI0/XI4/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_2 XI31/XI0/XI4/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI4/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_3 XI31/XI0/XI4/XI5/XI0/NET_0 XI31/XI0/XI4/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI4/XI5/XI0/MM_i_0 XI31/XI0/XI4/XI5/Z XI31/XI0/XI4/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI4/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI4/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI4/MUX0 XI31/XI0/XI4/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_6 XI31/XI0/XI4/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI4/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_9 XI31/XI0/XI4/XI5/XI0/NET_3 XI31/XI0/XI4/XI5/XI0/X1
+ XI31/XI0/XI4/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI4/MUX1 XI31/XI0/XI4/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI4/XI5/XI0/MM_i_1 XI31/XI0/XI4/XI5/Z XI31/XI0/XI4/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI4/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI4/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI4/XI3/MM_i_4 XI31/XI0/XI4/XI3/NET_1 XI31/XI0/XI4/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI3/MM_i_5 XI31/XI0/XI4/XI3/Z_NEG XI31/XI0/XI4/XI3/X1
+ XI31/XI0/XI4/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI3/MM_i_2 XI31/XI0/XI4/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI4/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI4/XI3/MM_i_3 XI31/XI0/XI4/XI3/NET_0 XI31/XI0/XI4/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI4/XI3/MM_i_0 XI31/XI0/XI4/MUX0 XI31/XI0/XI4/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI4/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI4/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI4/XI3/MM_i_8 VDD! XI31/XI0/XI4/NAND_OUT XI31/XI0/XI4/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI3/MM_i_6 XI31/XI0/XI4/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI4/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI3/MM_i_9 XI31/XI0/XI4/XI3/NET_3 XI31/XI0/XI4/XI3/X1
+ XI31/XI0/XI4/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI4/XI3/MM_i_7 VDD! XI31/XI0/XI4/XNOR_OUT XI31/XI0/XI4/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI4/XI3/MM_i_1 XI31/XI0/XI4/MUX0 XI31/XI0/XI4/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<1>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<14> ALU_OUT<1> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<1>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<14> ALU_OUT<1> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<1>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<14> ALU_OUT<1> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<1>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<14> ALU_OUT<1> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<1>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<14> ALU_OUT<1> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<1>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<14> ALU_OUT<1> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<1>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<14> ALU_OUT<1> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<1>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<14> ALU_OUT<1> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<1>/MM_i_0 XI31/XI2/NET3<14> XI31/XI2/ALU_PRE<1> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<1>/MM_i_1 XI31/XI2/NET3<14> XI31/XI2/ALU_PRE<1> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<1>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<1>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<1>/MM_i_4 XI31/XI2/XI0<1>/NET_1 XI31/LOGIC_OUT<1> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<1>/MM_i_5 XI31/XI2/XI0<1>/Z_NEG XI31/XI2/XI0<1>/X1
+ XI31/XI2/XI0<1>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<1>/MM_i_2 XI31/XI2/XI0<1>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<1>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<1>/MM_i_3 XI31/XI2/XI0<1>/NET_0 XI31/ARITHMETIC_OUT<1> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<1>/MM_i_0 XI31/XI2/ALU_PRE<1> XI31/XI2/XI0<1>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<1>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<1>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<1>/MM_i_8 VDD! XI31/LOGIC_OUT<1> XI31/XI2/XI0<1>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<1>/MM_i_6 XI31/XI2/XI0<1>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<1>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<1>/MM_i_9 XI31/XI2/XI0<1>/NET_3 XI31/XI2/XI0<1>/X1
+ XI31/XI2/XI0<1>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<1>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<1> XI31/XI2/XI0<1>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<1>/MM_i_1 XI31/XI2/ALU_PRE<1> XI31/XI2/XI0<1>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<0>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<15> ALU_OUT<0> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<0>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<15> ALU_OUT<0> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<0>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<15> ALU_OUT<0> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<0>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<15> ALU_OUT<0> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<0>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<15> ALU_OUT<0> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<0>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<15> ALU_OUT<0> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<0>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<15> ALU_OUT<0> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<0>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<15> ALU_OUT<0> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<0>/MM_i_0 XI31/XI2/NET3<15> XI31/XI2/ALU_PRE<0> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<0>/MM_i_1 XI31/XI2/NET3<15> XI31/XI2/ALU_PRE<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<0>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<0>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<0>/MM_i_4 XI31/XI2/XI0<0>/NET_1 XI31/LOGIC_OUT<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<0>/MM_i_5 XI31/XI2/XI0<0>/Z_NEG XI31/XI2/XI0<0>/X1
+ XI31/XI2/XI0<0>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<0>/MM_i_2 XI31/XI2/XI0<0>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<0>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<0>/MM_i_3 XI31/XI2/XI0<0>/NET_0 XI31/ARITHMETIC_OUT<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<0>/MM_i_0 XI31/XI2/ALU_PRE<0> XI31/XI2/XI0<0>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<0>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<0>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<0>/MM_i_8 VDD! XI31/LOGIC_OUT<0> XI31/XI2/XI0<0>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<0>/MM_i_6 XI31/XI2/XI0<0>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<0>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<0>/MM_i_9 XI31/XI2/XI0<0>/NET_3 XI31/XI2/XI0<0>/X1
+ XI31/XI2/XI0<0>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<0>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<0> XI31/XI2/XI0<0>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<0>/MM_i_1 XI31/XI2/ALU_PRE<0> XI31/XI2/XI0<0>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<3>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<12> ALU_OUT<3> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<3>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<12> ALU_OUT<3> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<3>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<12> ALU_OUT<3> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<3>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<12> ALU_OUT<3> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<3>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<12> ALU_OUT<3> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<3>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<12> ALU_OUT<3> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<3>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<12> ALU_OUT<3> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<3>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<12> ALU_OUT<3> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<3>/MM_i_0 XI31/XI2/NET3<12> XI31/XI2/ALU_PRE<3> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<3>/MM_i_1 XI31/XI2/NET3<12> XI31/XI2/ALU_PRE<3> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<3>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<3>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<3>/MM_i_4 XI31/XI2/XI0<3>/NET_1 XI31/LOGIC_OUT<3> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<3>/MM_i_5 XI31/XI2/XI0<3>/Z_NEG XI31/XI2/XI0<3>/X1
+ XI31/XI2/XI0<3>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<3>/MM_i_2 XI31/XI2/XI0<3>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<3>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<3>/MM_i_3 XI31/XI2/XI0<3>/NET_0 XI31/ARITHMETIC_OUT<3> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<3>/MM_i_0 XI31/XI2/ALU_PRE<3> XI31/XI2/XI0<3>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<3>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<3>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<3>/MM_i_8 VDD! XI31/LOGIC_OUT<3> XI31/XI2/XI0<3>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<3>/MM_i_6 XI31/XI2/XI0<3>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<3>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<3>/MM_i_9 XI31/XI2/XI0<3>/NET_3 XI31/XI2/XI0<3>/X1
+ XI31/XI2/XI0<3>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<3>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<3> XI31/XI2/XI0<3>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<3>/MM_i_1 XI31/XI2/ALU_PRE<3> XI31/XI2/XI0<3>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<2>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<13> ALU_OUT<2> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<2>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<13> ALU_OUT<2> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<2>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<13> ALU_OUT<2> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<2>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<13> ALU_OUT<2> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<2>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<13> ALU_OUT<2> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<2>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<13> ALU_OUT<2> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<2>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<13> ALU_OUT<2> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<2>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<13> ALU_OUT<2> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<2>/MM_i_0 XI31/XI2/NET3<13> XI31/XI2/ALU_PRE<2> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<2>/MM_i_1 XI31/XI2/NET3<13> XI31/XI2/ALU_PRE<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<2>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<2>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<2>/MM_i_4 XI31/XI2/XI0<2>/NET_1 XI31/LOGIC_OUT<2> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<2>/MM_i_5 XI31/XI2/XI0<2>/Z_NEG XI31/XI2/XI0<2>/X1
+ XI31/XI2/XI0<2>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<2>/MM_i_2 XI31/XI2/XI0<2>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<2>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<2>/MM_i_3 XI31/XI2/XI0<2>/NET_0 XI31/ARITHMETIC_OUT<2> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<2>/MM_i_0 XI31/XI2/ALU_PRE<2> XI31/XI2/XI0<2>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<2>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<2>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<2>/MM_i_8 VDD! XI31/LOGIC_OUT<2> XI31/XI2/XI0<2>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<2>/MM_i_6 XI31/XI2/XI0<2>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<2>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<2>/MM_i_9 XI31/XI2/XI0<2>/NET_3 XI31/XI2/XI0<2>/X1
+ XI31/XI2/XI0<2>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<2>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<2> XI31/XI2/XI0<2>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<2>/MM_i_1 XI31/XI2/ALU_PRE<2> XI31/XI2/XI0<2>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<5>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<10> ALU_OUT<5> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<5>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<10> ALU_OUT<5> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<5>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<10> ALU_OUT<5> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<5>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<10> ALU_OUT<5> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<5>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<10> ALU_OUT<5> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<5>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<10> ALU_OUT<5> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<5>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<10> ALU_OUT<5> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<5>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<10> ALU_OUT<5> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<5>/MM_i_0 XI31/XI2/NET3<10> XI31/XI2/ALU_PRE<5> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<5>/MM_i_1 XI31/XI2/NET3<10> XI31/XI2/ALU_PRE<5> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<5>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<5>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<5>/MM_i_4 XI31/XI2/XI0<5>/NET_1 XI31/LOGIC_OUT<5> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<5>/MM_i_5 XI31/XI2/XI0<5>/Z_NEG XI31/XI2/XI0<5>/X1
+ XI31/XI2/XI0<5>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<5>/MM_i_2 XI31/XI2/XI0<5>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<5>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<5>/MM_i_3 XI31/XI2/XI0<5>/NET_0 XI31/ARITHMETIC_OUT<5> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<5>/MM_i_0 XI31/XI2/ALU_PRE<5> XI31/XI2/XI0<5>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<5>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<5>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<5>/MM_i_8 VDD! XI31/LOGIC_OUT<5> XI31/XI2/XI0<5>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<5>/MM_i_6 XI31/XI2/XI0<5>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<5>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<5>/MM_i_9 XI31/XI2/XI0<5>/NET_3 XI31/XI2/XI0<5>/X1
+ XI31/XI2/XI0<5>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<5>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<5> XI31/XI2/XI0<5>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<5>/MM_i_1 XI31/XI2/ALU_PRE<5> XI31/XI2/XI0<5>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<4>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<11> ALU_OUT<4> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<4>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<11> ALU_OUT<4> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<4>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<11> ALU_OUT<4> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<4>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<11> ALU_OUT<4> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<4>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<11> ALU_OUT<4> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<4>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<11> ALU_OUT<4> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<4>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<11> ALU_OUT<4> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<4>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<11> ALU_OUT<4> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<4>/MM_i_0 XI31/XI2/NET3<11> XI31/XI2/ALU_PRE<4> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<4>/MM_i_1 XI31/XI2/NET3<11> XI31/XI2/ALU_PRE<4> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<4>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<4>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<4>/MM_i_4 XI31/XI2/XI0<4>/NET_1 XI31/LOGIC_OUT<4> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<4>/MM_i_5 XI31/XI2/XI0<4>/Z_NEG XI31/XI2/XI0<4>/X1
+ XI31/XI2/XI0<4>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<4>/MM_i_2 XI31/XI2/XI0<4>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<4>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<4>/MM_i_3 XI31/XI2/XI0<4>/NET_0 XI31/ARITHMETIC_OUT<4> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<4>/MM_i_0 XI31/XI2/ALU_PRE<4> XI31/XI2/XI0<4>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<4>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<4>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<4>/MM_i_8 VDD! XI31/LOGIC_OUT<4> XI31/XI2/XI0<4>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<4>/MM_i_6 XI31/XI2/XI0<4>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<4>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<4>/MM_i_9 XI31/XI2/XI0<4>/NET_3 XI31/XI2/XI0<4>/X1
+ XI31/XI2/XI0<4>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<4>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<4> XI31/XI2/XI0<4>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<4>/MM_i_1 XI31/XI2/ALU_PRE<4> XI31/XI2/XI0<4>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<7>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<8> ALU_OUT<7> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<7>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<8> ALU_OUT<7> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<7>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<8> ALU_OUT<7> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<7>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<8> ALU_OUT<7> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<7>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<8> ALU_OUT<7> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<7>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<8> ALU_OUT<7> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<7>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<8> ALU_OUT<7> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<7>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<8> ALU_OUT<7> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<7>/MM_i_0 XI31/XI2/NET3<8> XI31/XI2/ALU_PRE<7> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<7>/MM_i_1 XI31/XI2/NET3<8> XI31/XI2/ALU_PRE<7> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<7>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<7>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<7>/MM_i_4 XI31/XI2/XI0<7>/NET_1 XI31/LOGIC_OUT<7> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<7>/MM_i_5 XI31/XI2/XI0<7>/Z_NEG XI31/XI2/XI0<7>/X1
+ XI31/XI2/XI0<7>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<7>/MM_i_2 XI31/XI2/XI0<7>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<7>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<7>/MM_i_3 XI31/XI2/XI0<7>/NET_0 XI31/ARITHMETIC_OUT<7> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<7>/MM_i_0 XI31/XI2/ALU_PRE<7> XI31/XI2/XI0<7>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<7>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<7>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<7>/MM_i_8 VDD! XI31/LOGIC_OUT<7> XI31/XI2/XI0<7>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<7>/MM_i_6 XI31/XI2/XI0<7>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<7>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<7>/MM_i_9 XI31/XI2/XI0<7>/NET_3 XI31/XI2/XI0<7>/X1
+ XI31/XI2/XI0<7>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<7>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<7> XI31/XI2/XI0<7>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<7>/MM_i_1 XI31/XI2/ALU_PRE<7> XI31/XI2/XI0<7>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<6>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<9> ALU_OUT<6> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<6>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<9> ALU_OUT<6> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<6>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<9> ALU_OUT<6> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<6>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<9> ALU_OUT<6> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<6>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<9> ALU_OUT<6> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<6>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<9> ALU_OUT<6> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<6>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<9> ALU_OUT<6> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<6>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<9> ALU_OUT<6> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<6>/MM_i_0 XI31/XI2/NET3<9> XI31/XI2/ALU_PRE<6> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<6>/MM_i_1 XI31/XI2/NET3<9> XI31/XI2/ALU_PRE<6> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<6>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<6>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<6>/MM_i_4 XI31/XI2/XI0<6>/NET_1 XI31/LOGIC_OUT<6> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<6>/MM_i_5 XI31/XI2/XI0<6>/Z_NEG XI31/XI2/XI0<6>/X1
+ XI31/XI2/XI0<6>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<6>/MM_i_2 XI31/XI2/XI0<6>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<6>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<6>/MM_i_3 XI31/XI2/XI0<6>/NET_0 XI31/ARITHMETIC_OUT<6> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<6>/MM_i_0 XI31/XI2/ALU_PRE<6> XI31/XI2/XI0<6>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<6>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<6>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<6>/MM_i_8 VDD! XI31/LOGIC_OUT<6> XI31/XI2/XI0<6>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<6>/MM_i_6 XI31/XI2/XI0<6>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<6>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<6>/MM_i_9 XI31/XI2/XI0<6>/NET_3 XI31/XI2/XI0<6>/X1
+ XI31/XI2/XI0<6>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<6>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<6> XI31/XI2/XI0<6>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<6>/MM_i_1 XI31/XI2/ALU_PRE<6> XI31/XI2/XI0<6>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<9>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<6> ALU_OUT<9> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<9>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<6> ALU_OUT<9> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<9>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<6> ALU_OUT<9> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<9>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<6> ALU_OUT<9> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<9>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<6> ALU_OUT<9> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<9>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<6> ALU_OUT<9> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<9>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<6> ALU_OUT<9> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<9>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<6> ALU_OUT<9> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<9>/MM_i_0 XI31/XI2/NET3<6> XI31/XI2/ALU_PRE<9> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<9>/MM_i_1 XI31/XI2/NET3<6> XI31/XI2/ALU_PRE<9> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<9>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<9>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<9>/MM_i_4 XI31/XI2/XI0<9>/NET_1 XI31/LOGIC_OUT<9> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<9>/MM_i_5 XI31/XI2/XI0<9>/Z_NEG XI31/XI2/XI0<9>/X1
+ XI31/XI2/XI0<9>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<9>/MM_i_2 XI31/XI2/XI0<9>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<9>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<9>/MM_i_3 XI31/XI2/XI0<9>/NET_0 XI31/ARITHMETIC_OUT<9> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<9>/MM_i_0 XI31/XI2/ALU_PRE<9> XI31/XI2/XI0<9>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<9>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<9>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<9>/MM_i_8 VDD! XI31/LOGIC_OUT<9> XI31/XI2/XI0<9>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<9>/MM_i_6 XI31/XI2/XI0<9>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<9>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<9>/MM_i_9 XI31/XI2/XI0<9>/NET_3 XI31/XI2/XI0<9>/X1
+ XI31/XI2/XI0<9>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<9>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<9> XI31/XI2/XI0<9>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<9>/MM_i_1 XI31/XI2/ALU_PRE<9> XI31/XI2/XI0<9>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<8>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<7> ALU_OUT<8> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<8>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<7> ALU_OUT<8> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<8>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<7> ALU_OUT<8> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<8>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<7> ALU_OUT<8> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<8>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<7> ALU_OUT<8> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<8>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<7> ALU_OUT<8> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<8>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<7> ALU_OUT<8> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<8>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<7> ALU_OUT<8> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<8>/MM_i_0 XI31/XI2/NET3<7> XI31/XI2/ALU_PRE<8> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06
mXI31/XI2/XI1<8>/MM_i_1 XI31/XI2/NET3<7> XI31/XI2/ALU_PRE<8> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<8>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<8>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<8>/MM_i_4 XI31/XI2/XI0<8>/NET_1 XI31/LOGIC_OUT<8> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<8>/MM_i_5 XI31/XI2/XI0<8>/Z_NEG XI31/XI2/XI0<8>/X1
+ XI31/XI2/XI0<8>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<8>/MM_i_2 XI31/XI2/XI0<8>/Z_NEG CTRL_BUFF<2> XI31/XI2/XI0<8>/NET_0
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<8>/MM_i_3 XI31/XI2/XI0<8>/NET_0 XI31/ARITHMETIC_OUT<8> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<8>/MM_i_0 XI31/XI2/ALU_PRE<8> XI31/XI2/XI0<8>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<8>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<8>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<8>/MM_i_8 VDD! XI31/LOGIC_OUT<8> XI31/XI2/XI0<8>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<8>/MM_i_6 XI31/XI2/XI0<8>/NET_2 CTRL_BUFF<2> XI31/XI2/XI0<8>/Z_NEG
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<8>/MM_i_9 XI31/XI2/XI0<8>/NET_3 XI31/XI2/XI0<8>/X1
+ XI31/XI2/XI0<8>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14
+ PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<8>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<8> XI31/XI2/XI0<8>/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI2/XI0<8>/MM_i_1 XI31/XI2/ALU_PRE<8> XI31/XI2/XI0<8>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<11>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<4> ALU_OUT<11> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<11>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<4> ALU_OUT<11> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<11>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<4> ALU_OUT<11> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<11>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<4> ALU_OUT<11> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<11>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<4> ALU_OUT<11> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<11>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<4> ALU_OUT<11> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<11>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<4> ALU_OUT<11> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<11>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<4> ALU_OUT<11> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<11>/MM_i_0 XI31/XI2/NET3<4> XI31/XI2/ALU_PRE<11> VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI2/XI1<11>/MM_i_1 XI31/XI2/NET3<4> XI31/XI2/ALU_PRE<11> VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<11>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<11>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<11>/MM_i_4 XI31/XI2/XI0<11>/NET_1 XI31/LOGIC_OUT<11> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<11>/MM_i_5 XI31/XI2/XI0<11>/Z_NEG XI31/XI2/XI0<11>/X1
+ XI31/XI2/XI0<11>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<11>/MM_i_2 XI31/XI2/XI0<11>/Z_NEG CTRL_BUFF<2>
+ XI31/XI2/XI0<11>/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<11>/MM_i_3 XI31/XI2/XI0<11>/NET_0 XI31/ARITHMETIC_OUT<11> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<11>/MM_i_0 XI31/XI2/ALU_PRE<11> XI31/XI2/XI0<11>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<11>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<11>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<11>/MM_i_8 VDD! XI31/LOGIC_OUT<11> XI31/XI2/XI0<11>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<11>/MM_i_6 XI31/XI2/XI0<11>/NET_2 CTRL_BUFF<2>
+ XI31/XI2/XI0<11>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<11>/MM_i_9 XI31/XI2/XI0<11>/NET_3 XI31/XI2/XI0<11>/X1
+ XI31/XI2/XI0<11>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<11>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<11> XI31/XI2/XI0<11>/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI2/XI0<11>/MM_i_1 XI31/XI2/ALU_PRE<11> XI31/XI2/XI0<11>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<10>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<5> ALU_OUT<10> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<10>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<5> ALU_OUT<10> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<10>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<5> ALU_OUT<10> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<10>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<5> ALU_OUT<10> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<10>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<5> ALU_OUT<10> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<10>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<5> ALU_OUT<10> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<10>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<5> ALU_OUT<10> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<10>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<5> ALU_OUT<10> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<10>/MM_i_0 XI31/XI2/NET3<5> XI31/XI2/ALU_PRE<10> VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI2/XI1<10>/MM_i_1 XI31/XI2/NET3<5> XI31/XI2/ALU_PRE<10> VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<10>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<10>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<10>/MM_i_4 XI31/XI2/XI0<10>/NET_1 XI31/LOGIC_OUT<10> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<10>/MM_i_5 XI31/XI2/XI0<10>/Z_NEG XI31/XI2/XI0<10>/X1
+ XI31/XI2/XI0<10>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<10>/MM_i_2 XI31/XI2/XI0<10>/Z_NEG CTRL_BUFF<2>
+ XI31/XI2/XI0<10>/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<10>/MM_i_3 XI31/XI2/XI0<10>/NET_0 XI31/ARITHMETIC_OUT<10> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<10>/MM_i_0 XI31/XI2/ALU_PRE<10> XI31/XI2/XI0<10>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<10>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<10>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<10>/MM_i_8 VDD! XI31/LOGIC_OUT<10> XI31/XI2/XI0<10>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<10>/MM_i_6 XI31/XI2/XI0<10>/NET_2 CTRL_BUFF<2>
+ XI31/XI2/XI0<10>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<10>/MM_i_9 XI31/XI2/XI0<10>/NET_3 XI31/XI2/XI0<10>/X1
+ XI31/XI2/XI0<10>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<10>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<10> XI31/XI2/XI0<10>/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI2/XI0<10>/MM_i_1 XI31/XI2/ALU_PRE<10> XI31/XI2/XI0<10>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<13>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<2> ALU_OUT<13> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<13>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<2> ALU_OUT<13> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<13>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<2> ALU_OUT<13> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<13>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<2> ALU_OUT<13> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<13>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<2> ALU_OUT<13> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<13>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<2> ALU_OUT<13> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<13>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<2> ALU_OUT<13> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<13>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<2> ALU_OUT<13> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<13>/MM_i_0 XI31/XI2/NET3<2> XI31/XI2/ALU_PRE<13> VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI2/XI1<13>/MM_i_1 XI31/XI2/NET3<2> XI31/XI2/ALU_PRE<13> VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<13>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<13>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<13>/MM_i_4 XI31/XI2/XI0<13>/NET_1 XI31/LOGIC_OUT<13> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<13>/MM_i_5 XI31/XI2/XI0<13>/Z_NEG XI31/XI2/XI0<13>/X1
+ XI31/XI2/XI0<13>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<13>/MM_i_2 XI31/XI2/XI0<13>/Z_NEG CTRL_BUFF<2>
+ XI31/XI2/XI0<13>/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<13>/MM_i_3 XI31/XI2/XI0<13>/NET_0 XI31/ARITHMETIC_OUT<13> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<13>/MM_i_0 XI31/XI2/ALU_PRE<13> XI31/XI2/XI0<13>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<13>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<13>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<13>/MM_i_8 VDD! XI31/LOGIC_OUT<13> XI31/XI2/XI0<13>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<13>/MM_i_6 XI31/XI2/XI0<13>/NET_2 CTRL_BUFF<2>
+ XI31/XI2/XI0<13>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<13>/MM_i_9 XI31/XI2/XI0<13>/NET_3 XI31/XI2/XI0<13>/X1
+ XI31/XI2/XI0<13>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<13>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<13> XI31/XI2/XI0<13>/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI2/XI0<13>/MM_i_1 XI31/XI2/ALU_PRE<13> XI31/XI2/XI0<13>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<12>/MM_i_0_0_x4_0 VSS! XI31/XI2/NET3<3> ALU_OUT<12> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<12>/MM_i_0_0_x4_1 VSS! XI31/XI2/NET3<3> ALU_OUT<12> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<12>/MM_i_0_0_x4_2 VSS! XI31/XI2/NET3<3> ALU_OUT<12> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI2/XI2<12>/MM_i_0_0_x4_3 VSS! XI31/XI2/NET3<3> ALU_OUT<12> VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI2<12>/MM_i_1_0_x4_0 VDD! XI31/XI2/NET3<3> ALU_OUT<12> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI2<12>/MM_i_1_0_x4_1 VDD! XI31/XI2/NET3<3> ALU_OUT<12> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<12>/MM_i_1_0_x4_2 VDD! XI31/XI2/NET3<3> ALU_OUT<12> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI2/XI2<12>/MM_i_1_0_x4_3 VDD! XI31/XI2/NET3<3> ALU_OUT<12> VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI2/XI1<12>/MM_i_0 XI31/XI2/NET3<3> XI31/XI2/ALU_PRE<12> VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI2/XI1<12>/MM_i_1 XI31/XI2/NET3<3> XI31/XI2/ALU_PRE<12> VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI2/XI0<12>/MM_i_10 VSS! CTRL_BUFF<2> XI31/XI2/XI0<12>/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI2/XI0<12>/MM_i_4 XI31/XI2/XI0<12>/NET_1 XI31/LOGIC_OUT<12> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI2/XI0<12>/MM_i_5 XI31/XI2/XI0<12>/Z_NEG XI31/XI2/XI0<12>/X1
+ XI31/XI2/XI0<12>/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<12>/MM_i_2 XI31/XI2/XI0<12>/Z_NEG CTRL_BUFF<2>
+ XI31/XI2/XI0<12>/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI2/XI0<12>/MM_i_3 XI31/XI2/XI0<12>/NET_0 XI31/ARITHMETIC_OUT<12> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI2/XI0<12>/MM_i_0 XI31/XI2/ALU_PRE<12> XI31/XI2/XI0<12>/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI2/XI0<12>/MM_i_11 VDD! CTRL_BUFF<2> XI31/XI2/XI0<12>/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI2/XI0<12>/MM_i_8 VDD! XI31/LOGIC_OUT<12> XI31/XI2/XI0<12>/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<12>/MM_i_6 XI31/XI2/XI0<12>/NET_2 CTRL_BUFF<2>
+ XI31/XI2/XI0<12>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<12>/MM_i_9 XI31/XI2/XI0<12>/NET_3 XI31/XI2/XI0<12>/X1
+ XI31/XI2/XI0<12>/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI2/XI0<12>/MM_i_7 VDD! XI31/ARITHMETIC_OUT<12> XI31/XI2/XI0<12>/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI2/XI0<12>/MM_i_1 XI31/XI2/ALU_PRE<12> XI31/XI2/XI0<12>/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI15/XI0/MM_i_1 XI31/XI0/XI15/XI0/NET_0 OP0<0> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI15/XI0/MM_i_0 XI31/XI0/XI15/NAND_OUT OP1<0> XI31/XI0/XI15/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI15/XI1/MM_i_0 XI31/XI0/XI15/XI1/NET_001 OP1<0>
+ XI31/XI0/XI15/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI15/XI1/MM_i_5 VSS! OP0<0> XI31/XI0/XI15/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI15/XI1/MM_i_11 XI31/XI0/XI15/XI1/NET_002 XI31/XI0/XI15/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI15/XI1/MM_i_17 XI31/XI0/XI15/XNOR_OUT OP1<0>
+ XI31/XI0/XI15/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI15/XI1/MM_i_23 XI31/XI0/XI15/XI1/NET_002 OP0<0>
+ XI31/XI0/XI15/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI15/XI2/MM_i_1 XI31/XI0/XI15/NOR_OUT OP0<0> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI15/XI2/MM_i_0 VSS! OP1<0> XI31/XI0/XI15/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI15/XI0/MM_i_3 XI31/XI0/XI15/NAND_OUT OP0<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI15/XI0/MM_i_2 VDD! OP1<0> XI31/XI0/XI15/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI15/XI1/MM_i_29 XI31/XI0/XI15/XI1/NET_000 OP1<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI15/XI1/MM_i_36 VDD! OP0<0> XI31/XI0/XI15/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI15/XI1/MM_i_42 XI31/XI0/XI15/XNOR_OUT XI31/XI0/XI15/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI15/XI1/MM_i_48 XI31/XI0/XI15/XI1/NET_003 OP1<0>
+ XI31/XI0/XI15/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI15/XI1/MM_i_53 VDD! OP0<0> XI31/XI0/XI15/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI15/XI2/MM_i_3 XI31/XI0/XI15/XI2/NET_0 OP0<0> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI15/XI2/MM_i_2 XI31/XI0/XI15/NOR_OUT OP1<0> XI31/XI0/XI15/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI15/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<0> XI31/XI0/XI15/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI15/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<0> XI31/XI0/XI15/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI15/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI15/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI15/XI4/MM_i_4 XI31/XI0/XI15/XI4/NET_1 XI31/XI0/XI15/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI4/MM_i_5 XI31/XI0/XI15/XI4/Z_NEG XI31/XI0/XI15/XI4/X1
+ XI31/XI0/XI15/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI4/MM_i_2 XI31/XI0/XI15/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI15/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI4/MM_i_3 XI31/XI0/XI15/XI4/NET_0 OP0<0> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI15/XI4/MM_i_0 XI31/XI0/XI15/MUX1 XI31/XI0/XI15/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI15/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI15/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI15/XI4/MM_i_8 VDD! XI31/XI0/XI15/NOR_OUT XI31/XI0/XI15/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI4/MM_i_6 XI31/XI0/XI15/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI15/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI4/MM_i_9 XI31/XI0/XI15/XI4/NET_3 XI31/XI0/XI15/XI4/X1
+ XI31/XI0/XI15/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI4/MM_i_7 VDD! OP0<0> XI31/XI0/XI15/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI15/XI4/MM_i_1 XI31/XI0/XI15/MUX1 XI31/XI0/XI15/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI15/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI15/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_4 XI31/XI0/XI15/XI5/XI0/NET_1 XI31/XI0/XI15/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_5 XI31/XI0/XI15/XI5/XI0/Z_NEG
+ XI31/XI0/XI15/XI5/XI0/X1 XI31/XI0/XI15/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_2 XI31/XI0/XI15/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI15/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_3 XI31/XI0/XI15/XI5/XI0/NET_0 XI31/XI0/XI15/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI15/XI5/XI0/MM_i_0 XI31/XI0/XI15/XI5/Z XI31/XI0/XI15/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI15/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI15/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI15/MUX0
+ XI31/XI0/XI15/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_6 XI31/XI0/XI15/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI15/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_9 XI31/XI0/XI15/XI5/XI0/NET_3
+ XI31/XI0/XI15/XI5/XI0/X1 XI31/XI0/XI15/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI15/MUX1
+ XI31/XI0/XI15/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI15/XI5/XI0/MM_i_1 XI31/XI0/XI15/XI5/Z XI31/XI0/XI15/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI15/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI15/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI15/XI3/MM_i_4 XI31/XI0/XI15/XI3/NET_1 XI31/XI0/XI15/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI3/MM_i_5 XI31/XI0/XI15/XI3/Z_NEG XI31/XI0/XI15/XI3/X1
+ XI31/XI0/XI15/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI3/MM_i_2 XI31/XI0/XI15/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI15/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI15/XI3/MM_i_3 XI31/XI0/XI15/XI3/NET_0 XI31/XI0/XI15/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI15/XI3/MM_i_0 XI31/XI0/XI15/MUX0 XI31/XI0/XI15/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI15/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI15/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI15/XI3/MM_i_8 VDD! XI31/XI0/XI15/NAND_OUT XI31/XI0/XI15/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI3/MM_i_6 XI31/XI0/XI15/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI15/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI3/MM_i_9 XI31/XI0/XI15/XI3/NET_3 XI31/XI0/XI15/XI3/X1
+ XI31/XI0/XI15/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI15/XI3/MM_i_7 VDD! XI31/XI0/XI15/XNOR_OUT XI31/XI0/XI15/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI15/XI3/MM_i_1 XI31/XI0/XI15/MUX0 XI31/XI0/XI15/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI16/XI0/MM_i_1 XI31/XI0/XI16/XI0/NET_0 OP0<1> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI16/XI0/MM_i_0 XI31/XI0/XI16/NAND_OUT OP1<1> XI31/XI0/XI16/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI16/XI1/MM_i_0 XI31/XI0/XI16/XI1/NET_001 OP1<1>
+ XI31/XI0/XI16/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI16/XI1/MM_i_5 VSS! OP0<1> XI31/XI0/XI16/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI16/XI1/MM_i_11 XI31/XI0/XI16/XI1/NET_002 XI31/XI0/XI16/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI16/XI1/MM_i_17 XI31/XI0/XI16/XNOR_OUT OP1<1>
+ XI31/XI0/XI16/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI16/XI1/MM_i_23 XI31/XI0/XI16/XI1/NET_002 OP0<1>
+ XI31/XI0/XI16/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI16/XI2/MM_i_1 XI31/XI0/XI16/NOR_OUT OP0<1> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI16/XI2/MM_i_0 VSS! OP1<1> XI31/XI0/XI16/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI16/XI0/MM_i_3 XI31/XI0/XI16/NAND_OUT OP0<1> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI16/XI0/MM_i_2 VDD! OP1<1> XI31/XI0/XI16/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI16/XI1/MM_i_29 XI31/XI0/XI16/XI1/NET_000 OP1<1> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI16/XI1/MM_i_36 VDD! OP0<1> XI31/XI0/XI16/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI16/XI1/MM_i_42 XI31/XI0/XI16/XNOR_OUT XI31/XI0/XI16/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI16/XI1/MM_i_48 XI31/XI0/XI16/XI1/NET_003 OP1<1>
+ XI31/XI0/XI16/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI16/XI1/MM_i_53 VDD! OP0<1> XI31/XI0/XI16/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI16/XI2/MM_i_3 XI31/XI0/XI16/XI2/NET_0 OP0<1> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI16/XI2/MM_i_2 XI31/XI0/XI16/NOR_OUT OP1<1> XI31/XI0/XI16/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI16/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<1> XI31/XI0/XI16/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI16/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<1> XI31/XI0/XI16/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI16/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI16/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI16/XI4/MM_i_4 XI31/XI0/XI16/XI4/NET_1 XI31/XI0/XI16/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI4/MM_i_5 XI31/XI0/XI16/XI4/Z_NEG XI31/XI0/XI16/XI4/X1
+ XI31/XI0/XI16/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI4/MM_i_2 XI31/XI0/XI16/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI16/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI4/MM_i_3 XI31/XI0/XI16/XI4/NET_0 OP0<1> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI16/XI4/MM_i_0 XI31/XI0/XI16/MUX1 XI31/XI0/XI16/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI16/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI16/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI16/XI4/MM_i_8 VDD! XI31/XI0/XI16/NOR_OUT XI31/XI0/XI16/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI4/MM_i_6 XI31/XI0/XI16/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI16/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI4/MM_i_9 XI31/XI0/XI16/XI4/NET_3 XI31/XI0/XI16/XI4/X1
+ XI31/XI0/XI16/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI4/MM_i_7 VDD! OP0<1> XI31/XI0/XI16/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI16/XI4/MM_i_1 XI31/XI0/XI16/MUX1 XI31/XI0/XI16/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI16/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI16/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_4 XI31/XI0/XI16/XI5/XI0/NET_1 XI31/XI0/XI16/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_5 XI31/XI0/XI16/XI5/XI0/Z_NEG
+ XI31/XI0/XI16/XI5/XI0/X1 XI31/XI0/XI16/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_2 XI31/XI0/XI16/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI16/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_3 XI31/XI0/XI16/XI5/XI0/NET_0 XI31/XI0/XI16/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI16/XI5/XI0/MM_i_0 XI31/XI0/XI16/XI5/Z XI31/XI0/XI16/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI16/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI16/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI16/MUX0
+ XI31/XI0/XI16/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_6 XI31/XI0/XI16/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI16/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_9 XI31/XI0/XI16/XI5/XI0/NET_3
+ XI31/XI0/XI16/XI5/XI0/X1 XI31/XI0/XI16/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI16/MUX1
+ XI31/XI0/XI16/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI16/XI5/XI0/MM_i_1 XI31/XI0/XI16/XI5/Z XI31/XI0/XI16/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI16/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI16/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI16/XI3/MM_i_4 XI31/XI0/XI16/XI3/NET_1 XI31/XI0/XI16/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI3/MM_i_5 XI31/XI0/XI16/XI3/Z_NEG XI31/XI0/XI16/XI3/X1
+ XI31/XI0/XI16/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI3/MM_i_2 XI31/XI0/XI16/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI16/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI16/XI3/MM_i_3 XI31/XI0/XI16/XI3/NET_0 XI31/XI0/XI16/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI16/XI3/MM_i_0 XI31/XI0/XI16/MUX0 XI31/XI0/XI16/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI16/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI16/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI16/XI3/MM_i_8 VDD! XI31/XI0/XI16/NAND_OUT XI31/XI0/XI16/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI3/MM_i_6 XI31/XI0/XI16/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI16/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI3/MM_i_9 XI31/XI0/XI16/XI3/NET_3 XI31/XI0/XI16/XI3/X1
+ XI31/XI0/XI16/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI16/XI3/MM_i_7 VDD! XI31/XI0/XI16/XNOR_OUT XI31/XI0/XI16/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI16/XI3/MM_i_1 XI31/XI0/XI16/MUX0 XI31/XI0/XI16/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI14/XI0/MM_i_1 XI31/XI0/XI14/XI0/NET_0 OP0<2> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI14/XI0/MM_i_0 XI31/XI0/XI14/NAND_OUT OP1<2> XI31/XI0/XI14/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI14/XI1/MM_i_0 XI31/XI0/XI14/XI1/NET_001 OP1<2>
+ XI31/XI0/XI14/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI14/XI1/MM_i_5 VSS! OP0<2> XI31/XI0/XI14/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI14/XI1/MM_i_11 XI31/XI0/XI14/XI1/NET_002 XI31/XI0/XI14/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI14/XI1/MM_i_17 XI31/XI0/XI14/XNOR_OUT OP1<2>
+ XI31/XI0/XI14/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI14/XI1/MM_i_23 XI31/XI0/XI14/XI1/NET_002 OP0<2>
+ XI31/XI0/XI14/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI14/XI2/MM_i_1 XI31/XI0/XI14/NOR_OUT OP0<2> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI14/XI2/MM_i_0 VSS! OP1<2> XI31/XI0/XI14/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI14/XI0/MM_i_3 XI31/XI0/XI14/NAND_OUT OP0<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI14/XI0/MM_i_2 VDD! OP1<2> XI31/XI0/XI14/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI14/XI1/MM_i_29 XI31/XI0/XI14/XI1/NET_000 OP1<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI14/XI1/MM_i_36 VDD! OP0<2> XI31/XI0/XI14/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI14/XI1/MM_i_42 XI31/XI0/XI14/XNOR_OUT XI31/XI0/XI14/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI14/XI1/MM_i_48 XI31/XI0/XI14/XI1/NET_003 OP1<2>
+ XI31/XI0/XI14/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI14/XI1/MM_i_53 VDD! OP0<2> XI31/XI0/XI14/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI14/XI2/MM_i_3 XI31/XI0/XI14/XI2/NET_0 OP0<2> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI14/XI2/MM_i_2 XI31/XI0/XI14/NOR_OUT OP1<2> XI31/XI0/XI14/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI14/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<2> XI31/XI0/XI14/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI14/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<2> XI31/XI0/XI14/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI14/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI14/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI14/XI4/MM_i_4 XI31/XI0/XI14/XI4/NET_1 XI31/XI0/XI14/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI4/MM_i_5 XI31/XI0/XI14/XI4/Z_NEG XI31/XI0/XI14/XI4/X1
+ XI31/XI0/XI14/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI4/MM_i_2 XI31/XI0/XI14/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI14/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI4/MM_i_3 XI31/XI0/XI14/XI4/NET_0 OP0<2> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI14/XI4/MM_i_0 XI31/XI0/XI14/MUX1 XI31/XI0/XI14/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI14/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI14/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI14/XI4/MM_i_8 VDD! XI31/XI0/XI14/NOR_OUT XI31/XI0/XI14/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI4/MM_i_6 XI31/XI0/XI14/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI14/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI4/MM_i_9 XI31/XI0/XI14/XI4/NET_3 XI31/XI0/XI14/XI4/X1
+ XI31/XI0/XI14/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI4/MM_i_7 VDD! OP0<2> XI31/XI0/XI14/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI14/XI4/MM_i_1 XI31/XI0/XI14/MUX1 XI31/XI0/XI14/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI14/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI14/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_4 XI31/XI0/XI14/XI5/XI0/NET_1 XI31/XI0/XI14/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_5 XI31/XI0/XI14/XI5/XI0/Z_NEG
+ XI31/XI0/XI14/XI5/XI0/X1 XI31/XI0/XI14/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_2 XI31/XI0/XI14/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI14/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_3 XI31/XI0/XI14/XI5/XI0/NET_0 XI31/XI0/XI14/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI14/XI5/XI0/MM_i_0 XI31/XI0/XI14/XI5/Z XI31/XI0/XI14/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI14/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI14/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI14/MUX0
+ XI31/XI0/XI14/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_6 XI31/XI0/XI14/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI14/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_9 XI31/XI0/XI14/XI5/XI0/NET_3
+ XI31/XI0/XI14/XI5/XI0/X1 XI31/XI0/XI14/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI14/MUX1
+ XI31/XI0/XI14/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI14/XI5/XI0/MM_i_1 XI31/XI0/XI14/XI5/Z XI31/XI0/XI14/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI14/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI14/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI14/XI3/MM_i_4 XI31/XI0/XI14/XI3/NET_1 XI31/XI0/XI14/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI3/MM_i_5 XI31/XI0/XI14/XI3/Z_NEG XI31/XI0/XI14/XI3/X1
+ XI31/XI0/XI14/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI3/MM_i_2 XI31/XI0/XI14/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI14/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI14/XI3/MM_i_3 XI31/XI0/XI14/XI3/NET_0 XI31/XI0/XI14/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI14/XI3/MM_i_0 XI31/XI0/XI14/MUX0 XI31/XI0/XI14/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI14/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI14/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI14/XI3/MM_i_8 VDD! XI31/XI0/XI14/NAND_OUT XI31/XI0/XI14/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI3/MM_i_6 XI31/XI0/XI14/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI14/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI3/MM_i_9 XI31/XI0/XI14/XI3/NET_3 XI31/XI0/XI14/XI3/X1
+ XI31/XI0/XI14/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI14/XI3/MM_i_7 VDD! XI31/XI0/XI14/XNOR_OUT XI31/XI0/XI14/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI14/XI3/MM_i_1 XI31/XI0/XI14/MUX0 XI31/XI0/XI14/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI17/XI0/MM_i_1 XI31/XI0/XI17/XI0/NET_0 OP0<3> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI17/XI0/MM_i_0 XI31/XI0/XI17/NAND_OUT OP1<3> XI31/XI0/XI17/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI17/XI1/MM_i_0 XI31/XI0/XI17/XI1/NET_001 OP1<3>
+ XI31/XI0/XI17/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI17/XI1/MM_i_5 VSS! OP0<3> XI31/XI0/XI17/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI17/XI1/MM_i_11 XI31/XI0/XI17/XI1/NET_002 XI31/XI0/XI17/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI17/XI1/MM_i_17 XI31/XI0/XI17/XNOR_OUT OP1<3>
+ XI31/XI0/XI17/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI17/XI1/MM_i_23 XI31/XI0/XI17/XI1/NET_002 OP0<3>
+ XI31/XI0/XI17/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI17/XI2/MM_i_1 XI31/XI0/XI17/NOR_OUT OP0<3> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI17/XI2/MM_i_0 VSS! OP1<3> XI31/XI0/XI17/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI17/XI0/MM_i_3 XI31/XI0/XI17/NAND_OUT OP0<3> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI17/XI0/MM_i_2 VDD! OP1<3> XI31/XI0/XI17/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI17/XI1/MM_i_29 XI31/XI0/XI17/XI1/NET_000 OP1<3> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI17/XI1/MM_i_36 VDD! OP0<3> XI31/XI0/XI17/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI17/XI1/MM_i_42 XI31/XI0/XI17/XNOR_OUT XI31/XI0/XI17/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI17/XI1/MM_i_48 XI31/XI0/XI17/XI1/NET_003 OP1<3>
+ XI31/XI0/XI17/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI17/XI1/MM_i_53 VDD! OP0<3> XI31/XI0/XI17/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI17/XI2/MM_i_3 XI31/XI0/XI17/XI2/NET_0 OP0<3> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI17/XI2/MM_i_2 XI31/XI0/XI17/NOR_OUT OP1<3> XI31/XI0/XI17/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI17/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<3> XI31/XI0/XI17/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI17/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<3> XI31/XI0/XI17/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI17/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI17/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI17/XI4/MM_i_4 XI31/XI0/XI17/XI4/NET_1 XI31/XI0/XI17/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI4/MM_i_5 XI31/XI0/XI17/XI4/Z_NEG XI31/XI0/XI17/XI4/X1
+ XI31/XI0/XI17/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI4/MM_i_2 XI31/XI0/XI17/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI17/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI4/MM_i_3 XI31/XI0/XI17/XI4/NET_0 OP0<3> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI17/XI4/MM_i_0 XI31/XI0/XI17/MUX1 XI31/XI0/XI17/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI17/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI17/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI17/XI4/MM_i_8 VDD! XI31/XI0/XI17/NOR_OUT XI31/XI0/XI17/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI4/MM_i_6 XI31/XI0/XI17/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI17/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI4/MM_i_9 XI31/XI0/XI17/XI4/NET_3 XI31/XI0/XI17/XI4/X1
+ XI31/XI0/XI17/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI4/MM_i_7 VDD! OP0<3> XI31/XI0/XI17/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI17/XI4/MM_i_1 XI31/XI0/XI17/MUX1 XI31/XI0/XI17/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI17/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI17/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_4 XI31/XI0/XI17/XI5/XI0/NET_1 XI31/XI0/XI17/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_5 XI31/XI0/XI17/XI5/XI0/Z_NEG
+ XI31/XI0/XI17/XI5/XI0/X1 XI31/XI0/XI17/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_2 XI31/XI0/XI17/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI17/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_3 XI31/XI0/XI17/XI5/XI0/NET_0 XI31/XI0/XI17/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI17/XI5/XI0/MM_i_0 XI31/XI0/XI17/XI5/Z XI31/XI0/XI17/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI17/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI17/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI17/MUX0
+ XI31/XI0/XI17/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_6 XI31/XI0/XI17/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI17/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_9 XI31/XI0/XI17/XI5/XI0/NET_3
+ XI31/XI0/XI17/XI5/XI0/X1 XI31/XI0/XI17/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI17/MUX1
+ XI31/XI0/XI17/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI17/XI5/XI0/MM_i_1 XI31/XI0/XI17/XI5/Z XI31/XI0/XI17/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI17/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI17/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI17/XI3/MM_i_4 XI31/XI0/XI17/XI3/NET_1 XI31/XI0/XI17/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI3/MM_i_5 XI31/XI0/XI17/XI3/Z_NEG XI31/XI0/XI17/XI3/X1
+ XI31/XI0/XI17/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI3/MM_i_2 XI31/XI0/XI17/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI17/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI17/XI3/MM_i_3 XI31/XI0/XI17/XI3/NET_0 XI31/XI0/XI17/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI17/XI3/MM_i_0 XI31/XI0/XI17/MUX0 XI31/XI0/XI17/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI17/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI17/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI17/XI3/MM_i_8 VDD! XI31/XI0/XI17/NAND_OUT XI31/XI0/XI17/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI3/MM_i_6 XI31/XI0/XI17/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI17/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI3/MM_i_9 XI31/XI0/XI17/XI3/NET_3 XI31/XI0/XI17/XI3/X1
+ XI31/XI0/XI17/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI17/XI3/MM_i_7 VDD! XI31/XI0/XI17/XNOR_OUT XI31/XI0/XI17/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI17/XI3/MM_i_1 XI31/XI0/XI17/MUX0 XI31/XI0/XI17/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI12/XI0/MM_i_1 XI31/XI0/XI12/XI0/NET_0 OP0<4> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI12/XI0/MM_i_0 XI31/XI0/XI12/NAND_OUT OP1<4> XI31/XI0/XI12/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI12/XI1/MM_i_0 XI31/XI0/XI12/XI1/NET_001 OP1<4>
+ XI31/XI0/XI12/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI12/XI1/MM_i_5 VSS! OP0<4> XI31/XI0/XI12/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI12/XI1/MM_i_11 XI31/XI0/XI12/XI1/NET_002 XI31/XI0/XI12/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI12/XI1/MM_i_17 XI31/XI0/XI12/XNOR_OUT OP1<4>
+ XI31/XI0/XI12/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI12/XI1/MM_i_23 XI31/XI0/XI12/XI1/NET_002 OP0<4>
+ XI31/XI0/XI12/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI12/XI2/MM_i_1 XI31/XI0/XI12/NOR_OUT OP0<4> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI12/XI2/MM_i_0 VSS! OP1<4> XI31/XI0/XI12/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI12/XI0/MM_i_3 XI31/XI0/XI12/NAND_OUT OP0<4> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI12/XI0/MM_i_2 VDD! OP1<4> XI31/XI0/XI12/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI12/XI1/MM_i_29 XI31/XI0/XI12/XI1/NET_000 OP1<4> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI12/XI1/MM_i_36 VDD! OP0<4> XI31/XI0/XI12/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI12/XI1/MM_i_42 XI31/XI0/XI12/XNOR_OUT XI31/XI0/XI12/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI12/XI1/MM_i_48 XI31/XI0/XI12/XI1/NET_003 OP1<4>
+ XI31/XI0/XI12/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI12/XI1/MM_i_53 VDD! OP0<4> XI31/XI0/XI12/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI12/XI2/MM_i_3 XI31/XI0/XI12/XI2/NET_0 OP0<4> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI12/XI2/MM_i_2 XI31/XI0/XI12/NOR_OUT OP1<4> XI31/XI0/XI12/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI12/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<4> XI31/XI0/XI12/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI12/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<4> XI31/XI0/XI12/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI12/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI12/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI12/XI4/MM_i_4 XI31/XI0/XI12/XI4/NET_1 XI31/XI0/XI12/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI4/MM_i_5 XI31/XI0/XI12/XI4/Z_NEG XI31/XI0/XI12/XI4/X1
+ XI31/XI0/XI12/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI4/MM_i_2 XI31/XI0/XI12/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI12/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI4/MM_i_3 XI31/XI0/XI12/XI4/NET_0 OP0<4> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI12/XI4/MM_i_0 XI31/XI0/XI12/MUX1 XI31/XI0/XI12/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI12/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI12/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI12/XI4/MM_i_8 VDD! XI31/XI0/XI12/NOR_OUT XI31/XI0/XI12/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI4/MM_i_6 XI31/XI0/XI12/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI12/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI4/MM_i_9 XI31/XI0/XI12/XI4/NET_3 XI31/XI0/XI12/XI4/X1
+ XI31/XI0/XI12/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI4/MM_i_7 VDD! OP0<4> XI31/XI0/XI12/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI12/XI4/MM_i_1 XI31/XI0/XI12/MUX1 XI31/XI0/XI12/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI12/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI12/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_4 XI31/XI0/XI12/XI5/XI0/NET_1 XI31/XI0/XI12/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_5 XI31/XI0/XI12/XI5/XI0/Z_NEG
+ XI31/XI0/XI12/XI5/XI0/X1 XI31/XI0/XI12/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_2 XI31/XI0/XI12/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI12/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_3 XI31/XI0/XI12/XI5/XI0/NET_0 XI31/XI0/XI12/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI12/XI5/XI0/MM_i_0 XI31/XI0/XI12/XI5/Z XI31/XI0/XI12/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI12/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI12/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI12/MUX0
+ XI31/XI0/XI12/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_6 XI31/XI0/XI12/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI12/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_9 XI31/XI0/XI12/XI5/XI0/NET_3
+ XI31/XI0/XI12/XI5/XI0/X1 XI31/XI0/XI12/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI12/MUX1
+ XI31/XI0/XI12/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI12/XI5/XI0/MM_i_1 XI31/XI0/XI12/XI5/Z XI31/XI0/XI12/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI12/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI12/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI12/XI3/MM_i_4 XI31/XI0/XI12/XI3/NET_1 XI31/XI0/XI12/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI3/MM_i_5 XI31/XI0/XI12/XI3/Z_NEG XI31/XI0/XI12/XI3/X1
+ XI31/XI0/XI12/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI3/MM_i_2 XI31/XI0/XI12/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI12/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI12/XI3/MM_i_3 XI31/XI0/XI12/XI3/NET_0 XI31/XI0/XI12/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI12/XI3/MM_i_0 XI31/XI0/XI12/MUX0 XI31/XI0/XI12/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI12/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI12/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI12/XI3/MM_i_8 VDD! XI31/XI0/XI12/NAND_OUT XI31/XI0/XI12/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI3/MM_i_6 XI31/XI0/XI12/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI12/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI3/MM_i_9 XI31/XI0/XI12/XI3/NET_3 XI31/XI0/XI12/XI3/X1
+ XI31/XI0/XI12/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI12/XI3/MM_i_7 VDD! XI31/XI0/XI12/XNOR_OUT XI31/XI0/XI12/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI12/XI3/MM_i_1 XI31/XI0/XI12/MUX0 XI31/XI0/XI12/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI13/XI0/MM_i_1 XI31/XI0/XI13/XI0/NET_0 OP0<5> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI13/XI0/MM_i_0 XI31/XI0/XI13/NAND_OUT OP1<5> XI31/XI0/XI13/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI13/XI1/MM_i_0 XI31/XI0/XI13/XI1/NET_001 OP1<5>
+ XI31/XI0/XI13/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI13/XI1/MM_i_5 VSS! OP0<5> XI31/XI0/XI13/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI13/XI1/MM_i_11 XI31/XI0/XI13/XI1/NET_002 XI31/XI0/XI13/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI13/XI1/MM_i_17 XI31/XI0/XI13/XNOR_OUT OP1<5>
+ XI31/XI0/XI13/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI13/XI1/MM_i_23 XI31/XI0/XI13/XI1/NET_002 OP0<5>
+ XI31/XI0/XI13/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI13/XI2/MM_i_1 XI31/XI0/XI13/NOR_OUT OP0<5> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI13/XI2/MM_i_0 VSS! OP1<5> XI31/XI0/XI13/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI13/XI0/MM_i_3 XI31/XI0/XI13/NAND_OUT OP0<5> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI13/XI0/MM_i_2 VDD! OP1<5> XI31/XI0/XI13/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI13/XI1/MM_i_29 XI31/XI0/XI13/XI1/NET_000 OP1<5> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI13/XI1/MM_i_36 VDD! OP0<5> XI31/XI0/XI13/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI13/XI1/MM_i_42 XI31/XI0/XI13/XNOR_OUT XI31/XI0/XI13/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI13/XI1/MM_i_48 XI31/XI0/XI13/XI1/NET_003 OP1<5>
+ XI31/XI0/XI13/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI13/XI1/MM_i_53 VDD! OP0<5> XI31/XI0/XI13/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI13/XI2/MM_i_3 XI31/XI0/XI13/XI2/NET_0 OP0<5> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI13/XI2/MM_i_2 XI31/XI0/XI13/NOR_OUT OP1<5> XI31/XI0/XI13/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI13/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<5> XI31/XI0/XI13/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI13/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<5> XI31/XI0/XI13/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI13/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI13/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI13/XI4/MM_i_4 XI31/XI0/XI13/XI4/NET_1 XI31/XI0/XI13/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI4/MM_i_5 XI31/XI0/XI13/XI4/Z_NEG XI31/XI0/XI13/XI4/X1
+ XI31/XI0/XI13/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI4/MM_i_2 XI31/XI0/XI13/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI13/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI4/MM_i_3 XI31/XI0/XI13/XI4/NET_0 OP0<5> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI13/XI4/MM_i_0 XI31/XI0/XI13/MUX1 XI31/XI0/XI13/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI13/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI13/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI13/XI4/MM_i_8 VDD! XI31/XI0/XI13/NOR_OUT XI31/XI0/XI13/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI4/MM_i_6 XI31/XI0/XI13/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI13/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI4/MM_i_9 XI31/XI0/XI13/XI4/NET_3 XI31/XI0/XI13/XI4/X1
+ XI31/XI0/XI13/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI4/MM_i_7 VDD! OP0<5> XI31/XI0/XI13/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI13/XI4/MM_i_1 XI31/XI0/XI13/MUX1 XI31/XI0/XI13/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI13/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI13/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_4 XI31/XI0/XI13/XI5/XI0/NET_1 XI31/XI0/XI13/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_5 XI31/XI0/XI13/XI5/XI0/Z_NEG
+ XI31/XI0/XI13/XI5/XI0/X1 XI31/XI0/XI13/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_2 XI31/XI0/XI13/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI13/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_3 XI31/XI0/XI13/XI5/XI0/NET_0 XI31/XI0/XI13/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI13/XI5/XI0/MM_i_0 XI31/XI0/XI13/XI5/Z XI31/XI0/XI13/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI13/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI13/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI13/MUX0
+ XI31/XI0/XI13/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_6 XI31/XI0/XI13/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI13/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_9 XI31/XI0/XI13/XI5/XI0/NET_3
+ XI31/XI0/XI13/XI5/XI0/X1 XI31/XI0/XI13/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI13/MUX1
+ XI31/XI0/XI13/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI13/XI5/XI0/MM_i_1 XI31/XI0/XI13/XI5/Z XI31/XI0/XI13/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI13/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI13/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI13/XI3/MM_i_4 XI31/XI0/XI13/XI3/NET_1 XI31/XI0/XI13/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI3/MM_i_5 XI31/XI0/XI13/XI3/Z_NEG XI31/XI0/XI13/XI3/X1
+ XI31/XI0/XI13/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI3/MM_i_2 XI31/XI0/XI13/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI13/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI13/XI3/MM_i_3 XI31/XI0/XI13/XI3/NET_0 XI31/XI0/XI13/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI13/XI3/MM_i_0 XI31/XI0/XI13/MUX0 XI31/XI0/XI13/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI13/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI13/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI13/XI3/MM_i_8 VDD! XI31/XI0/XI13/NAND_OUT XI31/XI0/XI13/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI3/MM_i_6 XI31/XI0/XI13/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI13/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI3/MM_i_9 XI31/XI0/XI13/XI3/NET_3 XI31/XI0/XI13/XI3/X1
+ XI31/XI0/XI13/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI13/XI3/MM_i_7 VDD! XI31/XI0/XI13/XNOR_OUT XI31/XI0/XI13/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI13/XI3/MM_i_1 XI31/XI0/XI13/MUX0 XI31/XI0/XI13/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI11/XI0/MM_i_1 XI31/XI0/XI11/XI0/NET_0 OP0<6> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI11/XI0/MM_i_0 XI31/XI0/XI11/NAND_OUT OP1<6> XI31/XI0/XI11/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI11/XI1/MM_i_0 XI31/XI0/XI11/XI1/NET_001 OP1<6>
+ XI31/XI0/XI11/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI11/XI1/MM_i_5 VSS! OP0<6> XI31/XI0/XI11/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI11/XI1/MM_i_11 XI31/XI0/XI11/XI1/NET_002 XI31/XI0/XI11/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI11/XI1/MM_i_17 XI31/XI0/XI11/XNOR_OUT OP1<6>
+ XI31/XI0/XI11/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI11/XI1/MM_i_23 XI31/XI0/XI11/XI1/NET_002 OP0<6>
+ XI31/XI0/XI11/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI11/XI2/MM_i_1 XI31/XI0/XI11/NOR_OUT OP0<6> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI11/XI2/MM_i_0 VSS! OP1<6> XI31/XI0/XI11/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI11/XI0/MM_i_3 XI31/XI0/XI11/NAND_OUT OP0<6> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI11/XI0/MM_i_2 VDD! OP1<6> XI31/XI0/XI11/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI11/XI1/MM_i_29 XI31/XI0/XI11/XI1/NET_000 OP1<6> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI11/XI1/MM_i_36 VDD! OP0<6> XI31/XI0/XI11/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI11/XI1/MM_i_42 XI31/XI0/XI11/XNOR_OUT XI31/XI0/XI11/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI11/XI1/MM_i_48 XI31/XI0/XI11/XI1/NET_003 OP1<6>
+ XI31/XI0/XI11/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI11/XI1/MM_i_53 VDD! OP0<6> XI31/XI0/XI11/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI11/XI2/MM_i_3 XI31/XI0/XI11/XI2/NET_0 OP0<6> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI11/XI2/MM_i_2 XI31/XI0/XI11/NOR_OUT OP1<6> XI31/XI0/XI11/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI11/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<6> XI31/XI0/XI11/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI11/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<6> XI31/XI0/XI11/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI11/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI11/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI11/XI4/MM_i_4 XI31/XI0/XI11/XI4/NET_1 XI31/XI0/XI11/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI4/MM_i_5 XI31/XI0/XI11/XI4/Z_NEG XI31/XI0/XI11/XI4/X1
+ XI31/XI0/XI11/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI4/MM_i_2 XI31/XI0/XI11/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI11/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI4/MM_i_3 XI31/XI0/XI11/XI4/NET_0 OP0<6> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI11/XI4/MM_i_0 XI31/XI0/XI11/MUX1 XI31/XI0/XI11/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI11/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI11/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI11/XI4/MM_i_8 VDD! XI31/XI0/XI11/NOR_OUT XI31/XI0/XI11/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI4/MM_i_6 XI31/XI0/XI11/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI11/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI4/MM_i_9 XI31/XI0/XI11/XI4/NET_3 XI31/XI0/XI11/XI4/X1
+ XI31/XI0/XI11/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI4/MM_i_7 VDD! OP0<6> XI31/XI0/XI11/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI11/XI4/MM_i_1 XI31/XI0/XI11/MUX1 XI31/XI0/XI11/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI11/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI11/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_4 XI31/XI0/XI11/XI5/XI0/NET_1 XI31/XI0/XI11/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_5 XI31/XI0/XI11/XI5/XI0/Z_NEG
+ XI31/XI0/XI11/XI5/XI0/X1 XI31/XI0/XI11/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_2 XI31/XI0/XI11/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI11/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_3 XI31/XI0/XI11/XI5/XI0/NET_0 XI31/XI0/XI11/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI11/XI5/XI0/MM_i_0 XI31/XI0/XI11/XI5/Z XI31/XI0/XI11/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI11/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI11/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI11/MUX0
+ XI31/XI0/XI11/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_6 XI31/XI0/XI11/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI11/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_9 XI31/XI0/XI11/XI5/XI0/NET_3
+ XI31/XI0/XI11/XI5/XI0/X1 XI31/XI0/XI11/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI11/MUX1
+ XI31/XI0/XI11/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI11/XI5/XI0/MM_i_1 XI31/XI0/XI11/XI5/Z XI31/XI0/XI11/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI11/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI11/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI11/XI3/MM_i_4 XI31/XI0/XI11/XI3/NET_1 XI31/XI0/XI11/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI3/MM_i_5 XI31/XI0/XI11/XI3/Z_NEG XI31/XI0/XI11/XI3/X1
+ XI31/XI0/XI11/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI3/MM_i_2 XI31/XI0/XI11/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI11/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI11/XI3/MM_i_3 XI31/XI0/XI11/XI3/NET_0 XI31/XI0/XI11/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI11/XI3/MM_i_0 XI31/XI0/XI11/MUX0 XI31/XI0/XI11/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI11/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI11/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI11/XI3/MM_i_8 VDD! XI31/XI0/XI11/NAND_OUT XI31/XI0/XI11/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI3/MM_i_6 XI31/XI0/XI11/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI11/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI3/MM_i_9 XI31/XI0/XI11/XI3/NET_3 XI31/XI0/XI11/XI3/X1
+ XI31/XI0/XI11/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI11/XI3/MM_i_7 VDD! XI31/XI0/XI11/XNOR_OUT XI31/XI0/XI11/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI11/XI3/MM_i_1 XI31/XI0/XI11/MUX0 XI31/XI0/XI11/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI18/XI0/MM_i_1 XI31/XI0/XI18/XI0/NET_0 OP0<7> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI18/XI0/MM_i_0 XI31/XI0/XI18/NAND_OUT OP1<7> XI31/XI0/XI18/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI18/XI1/MM_i_0 XI31/XI0/XI18/XI1/NET_001 OP1<7>
+ XI31/XI0/XI18/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI18/XI1/MM_i_5 VSS! OP0<7> XI31/XI0/XI18/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI18/XI1/MM_i_11 XI31/XI0/XI18/XI1/NET_002 XI31/XI0/XI18/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI18/XI1/MM_i_17 XI31/XI0/XI18/XNOR_OUT OP1<7>
+ XI31/XI0/XI18/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI18/XI1/MM_i_23 XI31/XI0/XI18/XI1/NET_002 OP0<7>
+ XI31/XI0/XI18/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI18/XI2/MM_i_1 XI31/XI0/XI18/NOR_OUT OP0<7> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI18/XI2/MM_i_0 VSS! OP1<7> XI31/XI0/XI18/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI18/XI0/MM_i_3 XI31/XI0/XI18/NAND_OUT OP0<7> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI18/XI0/MM_i_2 VDD! OP1<7> XI31/XI0/XI18/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI18/XI1/MM_i_29 XI31/XI0/XI18/XI1/NET_000 OP1<7> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI18/XI1/MM_i_36 VDD! OP0<7> XI31/XI0/XI18/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI18/XI1/MM_i_42 XI31/XI0/XI18/XNOR_OUT XI31/XI0/XI18/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI18/XI1/MM_i_48 XI31/XI0/XI18/XI1/NET_003 OP1<7>
+ XI31/XI0/XI18/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI18/XI1/MM_i_53 VDD! OP0<7> XI31/XI0/XI18/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI18/XI2/MM_i_3 XI31/XI0/XI18/XI2/NET_0 OP0<7> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI18/XI2/MM_i_2 XI31/XI0/XI18/NOR_OUT OP1<7> XI31/XI0/XI18/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI18/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<7> XI31/XI0/XI18/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI18/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<7> XI31/XI0/XI18/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI18/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI18/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI18/XI4/MM_i_4 XI31/XI0/XI18/XI4/NET_1 XI31/XI0/XI18/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI4/MM_i_5 XI31/XI0/XI18/XI4/Z_NEG XI31/XI0/XI18/XI4/X1
+ XI31/XI0/XI18/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI4/MM_i_2 XI31/XI0/XI18/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI18/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI4/MM_i_3 XI31/XI0/XI18/XI4/NET_0 OP0<7> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI18/XI4/MM_i_0 XI31/XI0/XI18/MUX1 XI31/XI0/XI18/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI18/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI18/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI18/XI4/MM_i_8 VDD! XI31/XI0/XI18/NOR_OUT XI31/XI0/XI18/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI4/MM_i_6 XI31/XI0/XI18/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI18/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI4/MM_i_9 XI31/XI0/XI18/XI4/NET_3 XI31/XI0/XI18/XI4/X1
+ XI31/XI0/XI18/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI4/MM_i_7 VDD! OP0<7> XI31/XI0/XI18/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI18/XI4/MM_i_1 XI31/XI0/XI18/MUX1 XI31/XI0/XI18/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI18/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI18/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_4 XI31/XI0/XI18/XI5/XI0/NET_1 XI31/XI0/XI18/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_5 XI31/XI0/XI18/XI5/XI0/Z_NEG
+ XI31/XI0/XI18/XI5/XI0/X1 XI31/XI0/XI18/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_2 XI31/XI0/XI18/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI18/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_3 XI31/XI0/XI18/XI5/XI0/NET_0 XI31/XI0/XI18/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI18/XI5/XI0/MM_i_0 XI31/XI0/XI18/XI5/Z XI31/XI0/XI18/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI18/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI18/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI18/MUX0
+ XI31/XI0/XI18/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_6 XI31/XI0/XI18/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI18/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_9 XI31/XI0/XI18/XI5/XI0/NET_3
+ XI31/XI0/XI18/XI5/XI0/X1 XI31/XI0/XI18/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI18/MUX1
+ XI31/XI0/XI18/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI18/XI5/XI0/MM_i_1 XI31/XI0/XI18/XI5/Z XI31/XI0/XI18/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI18/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI18/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI18/XI3/MM_i_4 XI31/XI0/XI18/XI3/NET_1 XI31/XI0/XI18/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI3/MM_i_5 XI31/XI0/XI18/XI3/Z_NEG XI31/XI0/XI18/XI3/X1
+ XI31/XI0/XI18/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI3/MM_i_2 XI31/XI0/XI18/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI18/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI18/XI3/MM_i_3 XI31/XI0/XI18/XI3/NET_0 XI31/XI0/XI18/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI18/XI3/MM_i_0 XI31/XI0/XI18/MUX0 XI31/XI0/XI18/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI18/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI18/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI18/XI3/MM_i_8 VDD! XI31/XI0/XI18/NAND_OUT XI31/XI0/XI18/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI3/MM_i_6 XI31/XI0/XI18/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI18/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI3/MM_i_9 XI31/XI0/XI18/XI3/NET_3 XI31/XI0/XI18/XI3/X1
+ XI31/XI0/XI18/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI18/XI3/MM_i_7 VDD! XI31/XI0/XI18/XNOR_OUT XI31/XI0/XI18/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI18/XI3/MM_i_1 XI31/XI0/XI18/MUX0 XI31/XI0/XI18/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI8/XI0/MM_i_1 XI31/XI0/XI8/XI0/NET_0 OP0<8> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI8/XI0/MM_i_0 XI31/XI0/XI8/NAND_OUT OP1<8> XI31/XI0/XI8/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI8/XI1/MM_i_0 XI31/XI0/XI8/XI1/NET_001 OP1<8>
+ XI31/XI0/XI8/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI8/XI1/MM_i_5 VSS! OP0<8> XI31/XI0/XI8/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI8/XI1/MM_i_11 XI31/XI0/XI8/XI1/NET_002 XI31/XI0/XI8/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI8/XI1/MM_i_17 XI31/XI0/XI8/XNOR_OUT OP1<8> XI31/XI0/XI8/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI8/XI1/MM_i_23 XI31/XI0/XI8/XI1/NET_002 OP0<8> XI31/XI0/XI8/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI8/XI2/MM_i_1 XI31/XI0/XI8/NOR_OUT OP0<8> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI8/XI2/MM_i_0 VSS! OP1<8> XI31/XI0/XI8/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI8/XI0/MM_i_3 XI31/XI0/XI8/NAND_OUT OP0<8> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI8/XI0/MM_i_2 VDD! OP1<8> XI31/XI0/XI8/NAND_OUT VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI8/XI1/MM_i_29 XI31/XI0/XI8/XI1/NET_000 OP1<8> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI8/XI1/MM_i_36 VDD! OP0<8> XI31/XI0/XI8/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI8/XI1/MM_i_42 XI31/XI0/XI8/XNOR_OUT XI31/XI0/XI8/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI8/XI1/MM_i_48 XI31/XI0/XI8/XI1/NET_003 OP1<8> XI31/XI0/XI8/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI8/XI1/MM_i_53 VDD! OP0<8> XI31/XI0/XI8/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI8/XI2/MM_i_3 XI31/XI0/XI8/XI2/NET_0 OP0<8> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI8/XI2/MM_i_2 XI31/XI0/XI8/NOR_OUT OP1<8> XI31/XI0/XI8/XI2/NET_0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI8/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<8> XI31/XI0/XI8/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI8/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<8> XI31/XI0/XI8/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI8/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI8/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI8/XI4/MM_i_4 XI31/XI0/XI8/XI4/NET_1 XI31/XI0/XI8/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI4/MM_i_5 XI31/XI0/XI8/XI4/Z_NEG XI31/XI0/XI8/XI4/X1
+ XI31/XI0/XI8/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI4/MM_i_2 XI31/XI0/XI8/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI8/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI4/MM_i_3 XI31/XI0/XI8/XI4/NET_0 OP0<8> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI8/XI4/MM_i_0 XI31/XI0/XI8/MUX1 XI31/XI0/XI8/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI8/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI8/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI8/XI4/MM_i_8 VDD! XI31/XI0/XI8/NOR_OUT XI31/XI0/XI8/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI4/MM_i_6 XI31/XI0/XI8/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI8/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI4/MM_i_9 XI31/XI0/XI8/XI4/NET_3 XI31/XI0/XI8/XI4/X1
+ XI31/XI0/XI8/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI4/MM_i_7 VDD! OP0<8> XI31/XI0/XI8/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI8/XI4/MM_i_1 XI31/XI0/XI8/MUX1 XI31/XI0/XI8/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI8/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI8/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_4 XI31/XI0/XI8/XI5/XI0/NET_1 XI31/XI0/XI8/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_5 XI31/XI0/XI8/XI5/XI0/Z_NEG XI31/XI0/XI8/XI5/XI0/X1
+ XI31/XI0/XI8/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_2 XI31/XI0/XI8/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI8/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_3 XI31/XI0/XI8/XI5/XI0/NET_0 XI31/XI0/XI8/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI8/XI5/XI0/MM_i_0 XI31/XI0/XI8/XI5/Z XI31/XI0/XI8/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI8/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI8/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI8/MUX0 XI31/XI0/XI8/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_6 XI31/XI0/XI8/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI8/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_9 XI31/XI0/XI8/XI5/XI0/NET_3 XI31/XI0/XI8/XI5/XI0/X1
+ XI31/XI0/XI8/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI8/MUX1 XI31/XI0/XI8/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI8/XI5/XI0/MM_i_1 XI31/XI0/XI8/XI5/Z XI31/XI0/XI8/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI8/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI8/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI8/XI3/MM_i_4 XI31/XI0/XI8/XI3/NET_1 XI31/XI0/XI8/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI3/MM_i_5 XI31/XI0/XI8/XI3/Z_NEG XI31/XI0/XI8/XI3/X1
+ XI31/XI0/XI8/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI3/MM_i_2 XI31/XI0/XI8/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI8/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI8/XI3/MM_i_3 XI31/XI0/XI8/XI3/NET_0 XI31/XI0/XI8/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI8/XI3/MM_i_0 XI31/XI0/XI8/MUX0 XI31/XI0/XI8/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI8/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI8/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI8/XI3/MM_i_8 VDD! XI31/XI0/XI8/NAND_OUT XI31/XI0/XI8/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI3/MM_i_6 XI31/XI0/XI8/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI8/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI3/MM_i_9 XI31/XI0/XI8/XI3/NET_3 XI31/XI0/XI8/XI3/X1
+ XI31/XI0/XI8/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI8/XI3/MM_i_7 VDD! XI31/XI0/XI8/XNOR_OUT XI31/XI0/XI8/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI8/XI3/MM_i_1 XI31/XI0/XI8/MUX0 XI31/XI0/XI8/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI9/XI0/MM_i_1 XI31/XI0/XI9/XI0/NET_0 OP0<9> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI9/XI0/MM_i_0 XI31/XI0/XI9/NAND_OUT OP1<9> XI31/XI0/XI9/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI9/XI1/MM_i_0 XI31/XI0/XI9/XI1/NET_001 OP1<9>
+ XI31/XI0/XI9/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI9/XI1/MM_i_5 VSS! OP0<9> XI31/XI0/XI9/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI9/XI1/MM_i_11 XI31/XI0/XI9/XI1/NET_002 XI31/XI0/XI9/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI9/XI1/MM_i_17 XI31/XI0/XI9/XNOR_OUT OP1<9> XI31/XI0/XI9/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI9/XI1/MM_i_23 XI31/XI0/XI9/XI1/NET_002 OP0<9> XI31/XI0/XI9/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI9/XI2/MM_i_1 XI31/XI0/XI9/NOR_OUT OP0<9> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI9/XI2/MM_i_0 VSS! OP1<9> XI31/XI0/XI9/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI9/XI0/MM_i_3 XI31/XI0/XI9/NAND_OUT OP0<9> VDD! VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI9/XI0/MM_i_2 VDD! OP1<9> XI31/XI0/XI9/NAND_OUT VDD! PMOS_VTL L=5e-08
+ W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI9/XI1/MM_i_29 XI31/XI0/XI9/XI1/NET_000 OP1<9> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI9/XI1/MM_i_36 VDD! OP0<9> XI31/XI0/XI9/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI9/XI1/MM_i_42 XI31/XI0/XI9/XNOR_OUT XI31/XI0/XI9/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI9/XI1/MM_i_48 XI31/XI0/XI9/XI1/NET_003 OP1<9> XI31/XI0/XI9/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI9/XI1/MM_i_53 VDD! OP0<9> XI31/XI0/XI9/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI9/XI2/MM_i_3 XI31/XI0/XI9/XI2/NET_0 OP0<9> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI9/XI2/MM_i_2 XI31/XI0/XI9/NOR_OUT OP1<9> XI31/XI0/XI9/XI2/NET_0 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI9/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<9> XI31/XI0/XI9/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI9/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<9> XI31/XI0/XI9/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI9/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI9/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI9/XI4/MM_i_4 XI31/XI0/XI9/XI4/NET_1 XI31/XI0/XI9/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI4/MM_i_5 XI31/XI0/XI9/XI4/Z_NEG XI31/XI0/XI9/XI4/X1
+ XI31/XI0/XI9/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI4/MM_i_2 XI31/XI0/XI9/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI9/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI4/MM_i_3 XI31/XI0/XI9/XI4/NET_0 OP0<9> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI9/XI4/MM_i_0 XI31/XI0/XI9/MUX1 XI31/XI0/XI9/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI9/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI9/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI9/XI4/MM_i_8 VDD! XI31/XI0/XI9/NOR_OUT XI31/XI0/XI9/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI4/MM_i_6 XI31/XI0/XI9/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI9/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI4/MM_i_9 XI31/XI0/XI9/XI4/NET_3 XI31/XI0/XI9/XI4/X1
+ XI31/XI0/XI9/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI4/MM_i_7 VDD! OP0<9> XI31/XI0/XI9/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI9/XI4/MM_i_1 XI31/XI0/XI9/MUX1 XI31/XI0/XI9/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI9/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI9/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_4 XI31/XI0/XI9/XI5/XI0/NET_1 XI31/XI0/XI9/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_5 XI31/XI0/XI9/XI5/XI0/Z_NEG XI31/XI0/XI9/XI5/XI0/X1
+ XI31/XI0/XI9/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_2 XI31/XI0/XI9/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI9/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_3 XI31/XI0/XI9/XI5/XI0/NET_0 XI31/XI0/XI9/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI9/XI5/XI0/MM_i_0 XI31/XI0/XI9/XI5/Z XI31/XI0/XI9/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI9/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI9/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI9/MUX0 XI31/XI0/XI9/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_6 XI31/XI0/XI9/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI9/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_9 XI31/XI0/XI9/XI5/XI0/NET_3 XI31/XI0/XI9/XI5/XI0/X1
+ XI31/XI0/XI9/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI9/MUX1 XI31/XI0/XI9/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI9/XI5/XI0/MM_i_1 XI31/XI0/XI9/XI5/Z XI31/XI0/XI9/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI9/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI9/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI9/XI3/MM_i_4 XI31/XI0/XI9/XI3/NET_1 XI31/XI0/XI9/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI3/MM_i_5 XI31/XI0/XI9/XI3/Z_NEG XI31/XI0/XI9/XI3/X1
+ XI31/XI0/XI9/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI3/MM_i_2 XI31/XI0/XI9/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI9/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI9/XI3/MM_i_3 XI31/XI0/XI9/XI3/NET_0 XI31/XI0/XI9/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI9/XI3/MM_i_0 XI31/XI0/XI9/MUX0 XI31/XI0/XI9/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI9/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI9/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI9/XI3/MM_i_8 VDD! XI31/XI0/XI9/NAND_OUT XI31/XI0/XI9/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI3/MM_i_6 XI31/XI0/XI9/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI9/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI3/MM_i_9 XI31/XI0/XI9/XI3/NET_3 XI31/XI0/XI9/XI3/X1
+ XI31/XI0/XI9/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI9/XI3/MM_i_7 VDD! XI31/XI0/XI9/XNOR_OUT XI31/XI0/XI9/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI9/XI3/MM_i_1 XI31/XI0/XI9/MUX0 XI31/XI0/XI9/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI7/XI0/MM_i_1 XI31/XI0/XI7/XI0/NET_0 OP0<10> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI7/XI0/MM_i_0 XI31/XI0/XI7/NAND_OUT OP1<10> XI31/XI0/XI7/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI7/XI1/MM_i_0 XI31/XI0/XI7/XI1/NET_001 OP1<10>
+ XI31/XI0/XI7/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI7/XI1/MM_i_5 VSS! OP0<10> XI31/XI0/XI7/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI7/XI1/MM_i_11 XI31/XI0/XI7/XI1/NET_002 XI31/XI0/XI7/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI7/XI1/MM_i_17 XI31/XI0/XI7/XNOR_OUT OP1<10> XI31/XI0/XI7/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI7/XI1/MM_i_23 XI31/XI0/XI7/XI1/NET_002 OP0<10> XI31/XI0/XI7/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI7/XI2/MM_i_1 XI31/XI0/XI7/NOR_OUT OP0<10> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI7/XI2/MM_i_0 VSS! OP1<10> XI31/XI0/XI7/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI7/XI0/MM_i_3 XI31/XI0/XI7/NAND_OUT OP0<10> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI7/XI0/MM_i_2 VDD! OP1<10> XI31/XI0/XI7/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI7/XI1/MM_i_29 XI31/XI0/XI7/XI1/NET_000 OP1<10> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI7/XI1/MM_i_36 VDD! OP0<10> XI31/XI0/XI7/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI7/XI1/MM_i_42 XI31/XI0/XI7/XNOR_OUT XI31/XI0/XI7/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI7/XI1/MM_i_48 XI31/XI0/XI7/XI1/NET_003 OP1<10> XI31/XI0/XI7/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI7/XI1/MM_i_53 VDD! OP0<10> XI31/XI0/XI7/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI7/XI2/MM_i_3 XI31/XI0/XI7/XI2/NET_0 OP0<10> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI7/XI2/MM_i_2 XI31/XI0/XI7/NOR_OUT OP1<10> XI31/XI0/XI7/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI7/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<10> XI31/XI0/XI7/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI7/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<10> XI31/XI0/XI7/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI7/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI7/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI7/XI4/MM_i_4 XI31/XI0/XI7/XI4/NET_1 XI31/XI0/XI7/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI4/MM_i_5 XI31/XI0/XI7/XI4/Z_NEG XI31/XI0/XI7/XI4/X1
+ XI31/XI0/XI7/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI4/MM_i_2 XI31/XI0/XI7/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI7/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI4/MM_i_3 XI31/XI0/XI7/XI4/NET_0 OP0<10> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI7/XI4/MM_i_0 XI31/XI0/XI7/MUX1 XI31/XI0/XI7/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI7/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI7/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI7/XI4/MM_i_8 VDD! XI31/XI0/XI7/NOR_OUT XI31/XI0/XI7/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI4/MM_i_6 XI31/XI0/XI7/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI7/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI4/MM_i_9 XI31/XI0/XI7/XI4/NET_3 XI31/XI0/XI7/XI4/X1
+ XI31/XI0/XI7/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI4/MM_i_7 VDD! OP0<10> XI31/XI0/XI7/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI7/XI4/MM_i_1 XI31/XI0/XI7/MUX1 XI31/XI0/XI7/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI7/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI7/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_4 XI31/XI0/XI7/XI5/XI0/NET_1 XI31/XI0/XI7/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_5 XI31/XI0/XI7/XI5/XI0/Z_NEG XI31/XI0/XI7/XI5/XI0/X1
+ XI31/XI0/XI7/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_2 XI31/XI0/XI7/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI7/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_3 XI31/XI0/XI7/XI5/XI0/NET_0 XI31/XI0/XI7/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI7/XI5/XI0/MM_i_0 XI31/XI0/XI7/XI5/Z XI31/XI0/XI7/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI7/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI7/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI7/MUX0 XI31/XI0/XI7/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_6 XI31/XI0/XI7/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI7/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_9 XI31/XI0/XI7/XI5/XI0/NET_3 XI31/XI0/XI7/XI5/XI0/X1
+ XI31/XI0/XI7/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI7/MUX1 XI31/XI0/XI7/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI7/XI5/XI0/MM_i_1 XI31/XI0/XI7/XI5/Z XI31/XI0/XI7/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI7/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI7/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI7/XI3/MM_i_4 XI31/XI0/XI7/XI3/NET_1 XI31/XI0/XI7/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI3/MM_i_5 XI31/XI0/XI7/XI3/Z_NEG XI31/XI0/XI7/XI3/X1
+ XI31/XI0/XI7/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI3/MM_i_2 XI31/XI0/XI7/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI7/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI7/XI3/MM_i_3 XI31/XI0/XI7/XI3/NET_0 XI31/XI0/XI7/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI7/XI3/MM_i_0 XI31/XI0/XI7/MUX0 XI31/XI0/XI7/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI7/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI7/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI7/XI3/MM_i_8 VDD! XI31/XI0/XI7/NAND_OUT XI31/XI0/XI7/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI3/MM_i_6 XI31/XI0/XI7/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI7/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI3/MM_i_9 XI31/XI0/XI7/XI3/NET_3 XI31/XI0/XI7/XI3/X1
+ XI31/XI0/XI7/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI7/XI3/MM_i_7 VDD! XI31/XI0/XI7/XNOR_OUT XI31/XI0/XI7/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI7/XI3/MM_i_1 XI31/XI0/XI7/MUX0 XI31/XI0/XI7/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI10/XI0/MM_i_1 XI31/XI0/XI10/XI0/NET_0 OP0<11> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI10/XI0/MM_i_0 XI31/XI0/XI10/NAND_OUT OP1<11> XI31/XI0/XI10/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI10/XI1/MM_i_0 XI31/XI0/XI10/XI1/NET_001 OP1<11>
+ XI31/XI0/XI10/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI10/XI1/MM_i_5 VSS! OP0<11> XI31/XI0/XI10/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI10/XI1/MM_i_11 XI31/XI0/XI10/XI1/NET_002 XI31/XI0/XI10/XI1/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI10/XI1/MM_i_17 XI31/XI0/XI10/XNOR_OUT OP1<11>
+ XI31/XI0/XI10/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI0/XI10/XI1/MM_i_23 XI31/XI0/XI10/XI1/NET_002 OP0<11>
+ XI31/XI0/XI10/XNOR_OUT VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI10/XI2/MM_i_1 XI31/XI0/XI10/NOR_OUT OP0<11> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI10/XI2/MM_i_0 VSS! OP1<11> XI31/XI0/XI10/NOR_OUT VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI10/XI0/MM_i_3 XI31/XI0/XI10/NAND_OUT OP0<11> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI10/XI0/MM_i_2 VDD! OP1<11> XI31/XI0/XI10/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI10/XI1/MM_i_29 XI31/XI0/XI10/XI1/NET_000 OP1<11> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI10/XI1/MM_i_36 VDD! OP0<11> XI31/XI0/XI10/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI10/XI1/MM_i_42 XI31/XI0/XI10/XNOR_OUT XI31/XI0/XI10/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI10/XI1/MM_i_48 XI31/XI0/XI10/XI1/NET_003 OP1<11>
+ XI31/XI0/XI10/XNOR_OUT VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14
+ PD=1.54e-06 PS=1.54e-06
mXI31/XI0/XI10/XI1/MM_i_53 VDD! OP0<11> XI31/XI0/XI10/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI10/XI2/MM_i_3 XI31/XI0/XI10/XI2/NET_0 OP0<11> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI10/XI2/MM_i_2 XI31/XI0/XI10/NOR_OUT OP1<11> XI31/XI0/XI10/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI10/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<11> XI31/XI0/XI10/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI10/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<11> XI31/XI0/XI10/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI10/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI10/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI10/XI4/MM_i_4 XI31/XI0/XI10/XI4/NET_1 XI31/XI0/XI10/NOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI4/MM_i_5 XI31/XI0/XI10/XI4/Z_NEG XI31/XI0/XI10/XI4/X1
+ XI31/XI0/XI10/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI4/MM_i_2 XI31/XI0/XI10/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI10/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI4/MM_i_3 XI31/XI0/XI10/XI4/NET_0 OP0<11> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI10/XI4/MM_i_0 XI31/XI0/XI10/MUX1 XI31/XI0/XI10/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI10/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI10/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI10/XI4/MM_i_8 VDD! XI31/XI0/XI10/NOR_OUT XI31/XI0/XI10/XI4/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI4/MM_i_6 XI31/XI0/XI10/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI10/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI4/MM_i_9 XI31/XI0/XI10/XI4/NET_3 XI31/XI0/XI10/XI4/X1
+ XI31/XI0/XI10/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI4/MM_i_7 VDD! OP0<11> XI31/XI0/XI10/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI10/XI4/MM_i_1 XI31/XI0/XI10/MUX1 XI31/XI0/XI10/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI10/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI10/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_4 XI31/XI0/XI10/XI5/XI0/NET_1 XI31/XI0/XI10/MUX0
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_5 XI31/XI0/XI10/XI5/XI0/Z_NEG
+ XI31/XI0/XI10/XI5/XI0/X1 XI31/XI0/XI10/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_2 XI31/XI0/XI10/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI10/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_3 XI31/XI0/XI10/XI5/XI0/NET_0 XI31/XI0/XI10/MUX1
+ VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07
+ PS=1.11e-06
mXI31/XI0/XI10/XI5/XI0/MM_i_0 XI31/XI0/XI10/XI5/Z XI31/XI0/XI10/XI5/XI0/Z_NEG
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI10/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI10/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI10/MUX0
+ XI31/XI0/XI10/XI5/XI0/NET_2 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_6 XI31/XI0/XI10/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI10/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_9 XI31/XI0/XI10/XI5/XI0/NET_3
+ XI31/XI0/XI10/XI5/XI0/X1 XI31/XI0/XI10/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI10/MUX1
+ XI31/XI0/XI10/XI5/XI0/NET_3 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI10/XI5/XI0/MM_i_1 XI31/XI0/XI10/XI5/Z XI31/XI0/XI10/XI5/XI0/Z_NEG
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI10/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI10/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI10/XI3/MM_i_4 XI31/XI0/XI10/XI3/NET_1 XI31/XI0/XI10/NAND_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI3/MM_i_5 XI31/XI0/XI10/XI3/Z_NEG XI31/XI0/XI10/XI3/X1
+ XI31/XI0/XI10/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI3/MM_i_2 XI31/XI0/XI10/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI10/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI10/XI3/MM_i_3 XI31/XI0/XI10/XI3/NET_0 XI31/XI0/XI10/XNOR_OUT VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI10/XI3/MM_i_0 XI31/XI0/XI10/MUX0 XI31/XI0/XI10/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI10/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI10/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI10/XI3/MM_i_8 VDD! XI31/XI0/XI10/NAND_OUT XI31/XI0/XI10/XI3/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI3/MM_i_6 XI31/XI0/XI10/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI10/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI3/MM_i_9 XI31/XI0/XI10/XI3/NET_3 XI31/XI0/XI10/XI3/X1
+ XI31/XI0/XI10/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI10/XI3/MM_i_7 VDD! XI31/XI0/XI10/XNOR_OUT XI31/XI0/XI10/XI3/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI10/XI3/MM_i_1 XI31/XI0/XI10/MUX0 XI31/XI0/XI10/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI5/XI0/MM_i_1 XI31/XI0/XI5/XI0/NET_0 OP0<12> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI5/XI0/MM_i_0 XI31/XI0/XI5/NAND_OUT OP1<12> XI31/XI0/XI5/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI5/XI1/MM_i_0 XI31/XI0/XI5/XI1/NET_001 OP1<12>
+ XI31/XI0/XI5/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI5/XI1/MM_i_5 VSS! OP0<12> XI31/XI0/XI5/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI5/XI1/MM_i_11 XI31/XI0/XI5/XI1/NET_002 XI31/XI0/XI5/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI5/XI1/MM_i_17 XI31/XI0/XI5/XNOR_OUT OP1<12> XI31/XI0/XI5/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI5/XI1/MM_i_23 XI31/XI0/XI5/XI1/NET_002 OP0<12> XI31/XI0/XI5/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI5/XI2/MM_i_1 XI31/XI0/XI5/NOR_OUT OP0<12> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI5/XI2/MM_i_0 VSS! OP1<12> XI31/XI0/XI5/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI5/XI0/MM_i_3 XI31/XI0/XI5/NAND_OUT OP0<12> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI5/XI0/MM_i_2 VDD! OP1<12> XI31/XI0/XI5/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI5/XI1/MM_i_29 XI31/XI0/XI5/XI1/NET_000 OP1<12> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI5/XI1/MM_i_36 VDD! OP0<12> XI31/XI0/XI5/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI5/XI1/MM_i_42 XI31/XI0/XI5/XNOR_OUT XI31/XI0/XI5/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI5/XI1/MM_i_48 XI31/XI0/XI5/XI1/NET_003 OP1<12> XI31/XI0/XI5/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI5/XI1/MM_i_53 VDD! OP0<12> XI31/XI0/XI5/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI5/XI2/MM_i_3 XI31/XI0/XI5/XI2/NET_0 OP0<12> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI5/XI2/MM_i_2 XI31/XI0/XI5/NOR_OUT OP1<12> XI31/XI0/XI5/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI5/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<12> XI31/XI0/XI5/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI5/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<12> XI31/XI0/XI5/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI5/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI5/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI5/XI4/MM_i_4 XI31/XI0/XI5/XI4/NET_1 XI31/XI0/XI5/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI4/MM_i_5 XI31/XI0/XI5/XI4/Z_NEG XI31/XI0/XI5/XI4/X1
+ XI31/XI0/XI5/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI4/MM_i_2 XI31/XI0/XI5/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI5/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI4/MM_i_3 XI31/XI0/XI5/XI4/NET_0 OP0<12> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI5/XI4/MM_i_0 XI31/XI0/XI5/MUX1 XI31/XI0/XI5/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI5/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI5/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI5/XI4/MM_i_8 VDD! XI31/XI0/XI5/NOR_OUT XI31/XI0/XI5/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI4/MM_i_6 XI31/XI0/XI5/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI5/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI4/MM_i_9 XI31/XI0/XI5/XI4/NET_3 XI31/XI0/XI5/XI4/X1
+ XI31/XI0/XI5/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI4/MM_i_7 VDD! OP0<12> XI31/XI0/XI5/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI5/XI4/MM_i_1 XI31/XI0/XI5/MUX1 XI31/XI0/XI5/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI5/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI5/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_4 XI31/XI0/XI5/XI5/XI0/NET_1 XI31/XI0/XI5/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_5 XI31/XI0/XI5/XI5/XI0/Z_NEG XI31/XI0/XI5/XI5/XI0/X1
+ XI31/XI0/XI5/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_2 XI31/XI0/XI5/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI5/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_3 XI31/XI0/XI5/XI5/XI0/NET_0 XI31/XI0/XI5/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI5/XI5/XI0/MM_i_0 XI31/XI0/XI5/XI5/Z XI31/XI0/XI5/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI5/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI5/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI5/MUX0 XI31/XI0/XI5/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_6 XI31/XI0/XI5/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI5/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_9 XI31/XI0/XI5/XI5/XI0/NET_3 XI31/XI0/XI5/XI5/XI0/X1
+ XI31/XI0/XI5/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI5/MUX1 XI31/XI0/XI5/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI5/XI5/XI0/MM_i_1 XI31/XI0/XI5/XI5/Z XI31/XI0/XI5/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI5/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI5/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI5/XI3/MM_i_4 XI31/XI0/XI5/XI3/NET_1 XI31/XI0/XI5/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI3/MM_i_5 XI31/XI0/XI5/XI3/Z_NEG XI31/XI0/XI5/XI3/X1
+ XI31/XI0/XI5/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI3/MM_i_2 XI31/XI0/XI5/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI5/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI5/XI3/MM_i_3 XI31/XI0/XI5/XI3/NET_0 XI31/XI0/XI5/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI5/XI3/MM_i_0 XI31/XI0/XI5/MUX0 XI31/XI0/XI5/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI5/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI5/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI5/XI3/MM_i_8 VDD! XI31/XI0/XI5/NAND_OUT XI31/XI0/XI5/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI3/MM_i_6 XI31/XI0/XI5/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI5/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI3/MM_i_9 XI31/XI0/XI5/XI3/NET_3 XI31/XI0/XI5/XI3/X1
+ XI31/XI0/XI5/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI5/XI3/MM_i_7 VDD! XI31/XI0/XI5/XNOR_OUT XI31/XI0/XI5/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI5/XI3/MM_i_1 XI31/XI0/XI5/MUX0 XI31/XI0/XI5/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI6/XI0/MM_i_1 XI31/XI0/XI6/XI0/NET_0 OP0<13> VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI6/XI0/MM_i_0 XI31/XI0/XI6/NAND_OUT OP1<13> XI31/XI0/XI6/XI0/NET_0
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI6/XI1/MM_i_0 XI31/XI0/XI6/XI1/NET_001 OP1<13>
+ XI31/XI0/XI6/XI1/NET_000 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI6/XI1/MM_i_5 VSS! OP0<13> XI31/XI0/XI6/XI1/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI0/XI6/XI1/MM_i_11 XI31/XI0/XI6/XI1/NET_002 XI31/XI0/XI6/XI1/NET_000 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI0/XI6/XI1/MM_i_17 XI31/XI0/XI6/XNOR_OUT OP1<13> XI31/XI0/XI6/XI1/NET_002
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI0/XI6/XI1/MM_i_23 XI31/XI0/XI6/XI1/NET_002 OP0<13> XI31/XI0/XI6/XNOR_OUT
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI6/XI2/MM_i_1 XI31/XI0/XI6/NOR_OUT OP0<13> VSS! VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06
mXI31/XI0/XI6/XI2/MM_i_0 VSS! OP1<13> XI31/XI0/XI6/NOR_OUT VSS! NMOS_VTL L=5e-08
+ W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI6/XI0/MM_i_3 XI31/XI0/XI6/NAND_OUT OP0<13> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI6/XI0/MM_i_2 VDD! OP1<13> XI31/XI0/XI6/NAND_OUT VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI6/XI1/MM_i_29 XI31/XI0/XI6/XI1/NET_000 OP1<13> VDD! VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI6/XI1/MM_i_36 VDD! OP0<13> XI31/XI0/XI6/XI1/NET_000 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI0/XI6/XI1/MM_i_42 XI31/XI0/XI6/XNOR_OUT XI31/XI0/XI6/XI1/NET_000 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI0/XI6/XI1/MM_i_48 XI31/XI0/XI6/XI1/NET_003 OP1<13> XI31/XI0/XI6/XNOR_OUT
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI0/XI6/XI1/MM_i_53 VDD! OP0<13> XI31/XI0/XI6/XI1/NET_003 VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI6/XI2/MM_i_3 XI31/XI0/XI6/XI2/NET_0 OP0<13> VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06
mXI31/XI0/XI6/XI2/MM_i_2 XI31/XI0/XI6/NOR_OUT OP1<13> XI31/XI0/XI6/XI2/NET_0
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI6/XI5/XI1/MM_i_0 XI31/LOGIC_OUT<13> XI31/XI0/XI6/XI5/Z VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06
+ PS=1.04e-06
mXI31/XI0/XI6/XI5/XI1/MM_i_1 XI31/LOGIC_OUT<13> XI31/XI0/XI6/XI5/Z VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06
mXI31/XI0/XI6/XI4/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI6/XI4/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI6/XI4/MM_i_4 XI31/XI0/XI6/XI4/NET_1 XI31/XI0/XI6/NOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI4/MM_i_5 XI31/XI0/XI6/XI4/Z_NEG XI31/XI0/XI6/XI4/X1
+ XI31/XI0/XI6/XI4/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI4/MM_i_2 XI31/XI0/XI6/XI4/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI6/XI4/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI4/MM_i_3 XI31/XI0/XI6/XI4/NET_0 OP0<13> VSS! VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI6/XI4/MM_i_0 XI31/XI0/XI6/MUX1 XI31/XI0/XI6/XI4/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI6/XI4/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI6/XI4/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI6/XI4/MM_i_8 VDD! XI31/XI0/XI6/NOR_OUT XI31/XI0/XI6/XI4/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI4/MM_i_6 XI31/XI0/XI6/XI4/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI6/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI4/MM_i_9 XI31/XI0/XI6/XI4/NET_3 XI31/XI0/XI6/XI4/X1
+ XI31/XI0/XI6/XI4/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI4/MM_i_7 VDD! OP0<13> XI31/XI0/XI6/XI4/NET_3 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI6/XI4/MM_i_1 XI31/XI0/XI6/MUX1 XI31/XI0/XI6/XI4/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI0/XI6/XI5/XI0/MM_i_10 VSS! CTRL_BUFF<1> XI31/XI0/XI6/XI5/XI0/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_4 XI31/XI0/XI6/XI5/XI0/NET_1 XI31/XI0/XI6/MUX0 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_5 XI31/XI0/XI6/XI5/XI0/Z_NEG XI31/XI0/XI6/XI5/XI0/X1
+ XI31/XI0/XI6/XI5/XI0/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_2 XI31/XI0/XI6/XI5/XI0/Z_NEG CTRL_BUFF<1>
+ XI31/XI0/XI6/XI5/XI0/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_3 XI31/XI0/XI6/XI5/XI0/NET_0 XI31/XI0/XI6/MUX1 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI6/XI5/XI0/MM_i_0 XI31/XI0/XI6/XI5/Z XI31/XI0/XI6/XI5/XI0/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI0/XI6/XI5/XI0/MM_i_11 VDD! CTRL_BUFF<1> XI31/XI0/XI6/XI5/XI0/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_8 VDD! XI31/XI0/XI6/MUX0 XI31/XI0/XI6/XI5/XI0/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_6 XI31/XI0/XI6/XI5/XI0/NET_2 CTRL_BUFF<1>
+ XI31/XI0/XI6/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_9 XI31/XI0/XI6/XI5/XI0/NET_3 XI31/XI0/XI6/XI5/XI0/X1
+ XI31/XI0/XI6/XI5/XI0/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_7 VDD! XI31/XI0/XI6/MUX1 XI31/XI0/XI6/XI5/XI0/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI0/XI6/XI5/XI0/MM_i_1 XI31/XI0/XI6/XI5/Z XI31/XI0/XI6/XI5/XI0/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI0/XI6/XI3/MM_i_10 VSS! CTRL_BUFF<0> XI31/XI0/XI6/XI3/X1 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI0/XI6/XI3/MM_i_4 XI31/XI0/XI6/XI3/NET_1 XI31/XI0/XI6/NAND_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI3/MM_i_5 XI31/XI0/XI6/XI3/Z_NEG XI31/XI0/XI6/XI3/X1
+ XI31/XI0/XI6/XI3/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI3/MM_i_2 XI31/XI0/XI6/XI3/Z_NEG CTRL_BUFF<0>
+ XI31/XI0/XI6/XI3/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14
+ PD=7e-07 PS=7e-07
mXI31/XI0/XI6/XI3/MM_i_3 XI31/XI0/XI6/XI3/NET_0 XI31/XI0/XI6/XNOR_OUT VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI0/XI6/XI3/MM_i_0 XI31/XI0/XI6/MUX0 XI31/XI0/XI6/XI3/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI0/XI6/XI3/MM_i_11 VDD! CTRL_BUFF<0> XI31/XI0/XI6/XI3/X1 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI0/XI6/XI3/MM_i_8 VDD! XI31/XI0/XI6/NAND_OUT XI31/XI0/XI6/XI3/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI3/MM_i_6 XI31/XI0/XI6/XI3/NET_2 CTRL_BUFF<0>
+ XI31/XI0/XI6/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI3/MM_i_9 XI31/XI0/XI6/XI3/NET_3 XI31/XI0/XI6/XI3/X1
+ XI31/XI0/XI6/XI3/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI0/XI6/XI3/MM_i_7 VDD! XI31/XI0/XI6/XNOR_OUT XI31/XI0/XI6/XI3/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI0/XI6/XI3/MM_i_1 XI31/XI0/XI6/MUX0 XI31/XI0/XI6/XI3/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI40/XI9/MM_i_0 XI31/XI1/XI40/XI9/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI40/XI9/MM_i_7 VSS! OP0<0> XI31/XI1/XI40/XI9/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI40/XI9/MM_i_13 XI31/XI1/XI40/OP0_TEMP<0> XI31/XI1/XI40/XI9/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI40/XI9/MM_i_19 XI31/XI1/XI40/XI9/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI40/OP0_TEMP<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI40/XI9/MM_i_24 VSS! OP0<0> XI31/XI1/XI40/XI9/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI40/XI9/MM_i_30 XI31/XI1/XI40/XI9/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI40/XI9/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI40/XI9/MM_i_35 VDD! OP0<0> XI31/XI1/XI40/XI9/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI40/XI9/MM_i_41 XI31/XI1/XI40/XI9/NET_003 XI31/XI1/XI40/XI9/NET_000
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI1/XI40/XI9/MM_i_47 XI31/XI1/XI40/OP0_TEMP<0> CTRL_BUFF<0>
+ XI31/XI1/XI40/XI9/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI40/XI9/MM_i_53 XI31/XI1/XI40/XI9/NET_003 OP0<0>
+ XI31/XI1/XI40/OP0_TEMP<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI40/XI10/MM_i_0 XI31/XI1/XI40/XI10/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI40/XI10/MM_i_7 VSS! OP0<1> XI31/XI1/XI40/XI10/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI40/XI10/MM_i_13 XI31/XI1/XI40/OP0_TEMP<1> XI31/XI1/XI40/XI10/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI40/XI10/MM_i_19 XI31/XI1/XI40/XI10/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI40/OP0_TEMP<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI40/XI10/MM_i_24 VSS! OP0<1> XI31/XI1/XI40/XI10/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI40/XI10/MM_i_30 XI31/XI1/XI40/XI10/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI40/XI10/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI40/XI10/MM_i_35 VDD! OP0<1> XI31/XI1/XI40/XI10/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI40/XI10/MM_i_41 XI31/XI1/XI40/XI10/NET_003
+ XI31/XI1/XI40/XI10/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI40/XI10/MM_i_47 XI31/XI1/XI40/OP0_TEMP<1> CTRL_BUFF<0>
+ XI31/XI1/XI40/XI10/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI40/XI10/MM_i_53 XI31/XI1/XI40/XI10/NET_003 OP0<1>
+ XI31/XI1/XI40/OP0_TEMP<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI40/XI0/MM_instance_159 XI31/XI1/XI40/NET16 XI31/XI1/XI40/XI0/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI40/XI0/MM_instance_166 VSS! OP1<0> XI31/XI1/XI40/XI0/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_170 XI31/XI1/XI40/XI0/NET_000
+ XI31/XI1/XI40/OP0_TEMP<0> XI31/XI1/XI40/XI0/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_176 XI31/XI1/XI40/XI0/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI40/XI0/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI40/XI0/MM_instance_188 XI31/XI1/XI40/XI0/NET_002
+ XI31/XI1/XI40/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_182 VSS! OP1<0> XI31/XI1/XI40/XI0/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI40/XI0/MM_instance_227 XI31/XI1/XI40/XI0/NET_006 OP1<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI40/XI0/MM_instance_215 VSS! CTRL_BUFF<0> XI31/XI1/XI40/XI0/NET_006
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_221 XI31/XI1/XI40/XI0/NET_006
+ XI31/XI1/XI40/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_209 XI31/XI1/XI40/XI0/NET_005
+ XI31/XI1/XI40/XI0/NET_001 XI31/XI1/XI40/XI0/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_203 XI31/XI1/XI40/XI0/NET_004 CTRL_BUFF<0>
+ XI31/XI1/XI40/XI0/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI40/XI0/MM_instance_199 XI31/XI1/XI40/XI0/NET_003 OP1<0>
+ XI31/XI1/XI40/XI0/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_194 VSS! XI31/XI1/XI40/OP0_TEMP<0>
+ XI31/XI1/XI40/XI0/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI40/XI0/MM_instance_233 XI31/ARITHMETIC_OUT<0>
+ XI31/XI1/XI40/XI0/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI40/XI0/MM_instance_239 XI31/XI1/XI40/NET16 XI31/XI1/XI40/XI0/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI40/XI0/MM_instance_246 VDD! OP1<0> XI31/XI1/XI40/XI0/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_251 XI31/XI1/XI40/XI0/NET_007
+ XI31/XI1/XI40/OP0_TEMP<0> XI31/XI1/XI40/XI0/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_257 XI31/XI1/XI40/XI0/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI40/XI0/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI40/XI0/MM_instance_269 XI31/XI1/XI40/XI0/NET_008
+ XI31/XI1/XI40/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_263 VDD! OP1<0> XI31/XI1/XI40/XI0/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI40/XI0/MM_instance_309 XI31/XI1/XI40/XI0/NET_011 OP1<0> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI40/XI0/MM_instance_297 VDD! CTRL_BUFF<0> XI31/XI1/XI40/XI0/NET_011
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_303 XI31/XI1/XI40/XI0/NET_011
+ XI31/XI1/XI40/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_290 XI31/XI1/XI40/XI0/NET_005
+ XI31/XI1/XI40/XI0/NET_001 XI31/XI1/XI40/XI0/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_284 XI31/XI1/XI40/XI0/NET_010 CTRL_BUFF<0>
+ XI31/XI1/XI40/XI0/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI40/XI0/MM_instance_280 XI31/XI1/XI40/XI0/NET_009 OP1<0>
+ XI31/XI1/XI40/XI0/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_275 VDD! XI31/XI1/XI40/OP0_TEMP<0>
+ XI31/XI1/XI40/XI0/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI40/XI0/MM_instance_315 XI31/ARITHMETIC_OUT<0>
+ XI31/XI1/XI40/XI0/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI40/XI1/MM_instance_159 XI31/XI1/NET1 XI31/XI1/XI40/XI1/NET_001 VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI40/XI1/MM_instance_166 VSS! OP1<1> XI31/XI1/XI40/XI1/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_170 XI31/XI1/XI40/XI1/NET_000
+ XI31/XI1/XI40/OP0_TEMP<1> XI31/XI1/XI40/XI1/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_176 XI31/XI1/XI40/XI1/NET_001 XI31/XI1/XI40/NET16
+ XI31/XI1/XI40/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI40/XI1/MM_instance_188 XI31/XI1/XI40/XI1/NET_002
+ XI31/XI1/XI40/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_182 VSS! OP1<1> XI31/XI1/XI40/XI1/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI40/XI1/MM_instance_227 XI31/XI1/XI40/XI1/NET_006 OP1<1> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI40/XI1/MM_instance_215 VSS! XI31/XI1/XI40/NET16
+ XI31/XI1/XI40/XI1/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_221 XI31/XI1/XI40/XI1/NET_006
+ XI31/XI1/XI40/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_209 XI31/XI1/XI40/XI1/NET_005
+ XI31/XI1/XI40/XI1/NET_001 XI31/XI1/XI40/XI1/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_203 XI31/XI1/XI40/XI1/NET_004 XI31/XI1/XI40/NET16
+ XI31/XI1/XI40/XI1/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI40/XI1/MM_instance_199 XI31/XI1/XI40/XI1/NET_003 OP1<1>
+ XI31/XI1/XI40/XI1/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_194 VSS! XI31/XI1/XI40/OP0_TEMP<1>
+ XI31/XI1/XI40/XI1/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI40/XI1/MM_instance_233 XI31/ARITHMETIC_OUT<1>
+ XI31/XI1/XI40/XI1/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI40/XI1/MM_instance_239 XI31/XI1/NET1 XI31/XI1/XI40/XI1/NET_001 VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI40/XI1/MM_instance_246 VDD! OP1<1> XI31/XI1/XI40/XI1/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_251 XI31/XI1/XI40/XI1/NET_007
+ XI31/XI1/XI40/OP0_TEMP<1> XI31/XI1/XI40/XI1/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_257 XI31/XI1/XI40/XI1/NET_001 XI31/XI1/XI40/NET16
+ XI31/XI1/XI40/XI1/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI40/XI1/MM_instance_269 XI31/XI1/XI40/XI1/NET_008
+ XI31/XI1/XI40/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_263 VDD! OP1<1> XI31/XI1/XI40/XI1/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI40/XI1/MM_instance_309 XI31/XI1/XI40/XI1/NET_011 OP1<1> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI40/XI1/MM_instance_297 VDD! XI31/XI1/XI40/NET16
+ XI31/XI1/XI40/XI1/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_303 XI31/XI1/XI40/XI1/NET_011
+ XI31/XI1/XI40/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_290 XI31/XI1/XI40/XI1/NET_005
+ XI31/XI1/XI40/XI1/NET_001 XI31/XI1/XI40/XI1/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_284 XI31/XI1/XI40/XI1/NET_010 XI31/XI1/XI40/NET16
+ XI31/XI1/XI40/XI1/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI40/XI1/MM_instance_280 XI31/XI1/XI40/XI1/NET_009 OP1<1>
+ XI31/XI1/XI40/XI1/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_275 VDD! XI31/XI1/XI40/OP0_TEMP<1>
+ XI31/XI1/XI40/XI1/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI40/XI1/MM_instance_315 XI31/ARITHMETIC_OUT<1>
+ XI31/XI1/XI40/XI1/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI17/MM_i_10 VSS! XI31/XI1/NET16 XI31/XI1/XI44/XI17/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI17/MM_i_4 XI31/XI1/XI44/XI17/NET_1 XI31/XI1/XI44/S_0<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI17/MM_i_5 XI31/XI1/XI44/XI17/Z_NEG XI31/XI1/XI44/XI17/X1
+ XI31/XI1/XI44/XI17/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI17/MM_i_2 XI31/XI1/XI44/XI17/Z_NEG XI31/XI1/NET16
+ XI31/XI1/XI44/XI17/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI17/MM_i_3 XI31/XI1/XI44/XI17/NET_0 XI31/XI1/XI44/S_1<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI44/XI17/MM_i_0 XI31/ARITHMETIC_OUT<11> XI31/XI1/XI44/XI17/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI17/MM_i_11 VDD! XI31/XI1/NET16 XI31/XI1/XI44/XI17/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI17/MM_i_8 VDD! XI31/XI1/XI44/S_0<0> XI31/XI1/XI44/XI17/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI17/MM_i_6 XI31/XI1/XI44/XI17/NET_2 XI31/XI1/NET16
+ XI31/XI1/XI44/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI17/MM_i_9 XI31/XI1/XI44/XI17/NET_3 XI31/XI1/XI44/XI17/X1
+ XI31/XI1/XI44/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI17/MM_i_7 VDD! XI31/XI1/XI44/S_1<0> XI31/XI1/XI44/XI17/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI17/MM_i_1 XI31/ARITHMETIC_OUT<11> XI31/XI1/XI44/XI17/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI25/MM_i_10 VSS! XI31/XI1/NET16 XI31/XI1/XI44/XI25/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI25/MM_i_4 XI31/XI1/XI44/XI25/NET_1 XI31/XI1/XI44/S_0<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI25/MM_i_5 XI31/XI1/XI44/XI25/Z_NEG XI31/XI1/XI44/XI25/X1
+ XI31/XI1/XI44/XI25/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI25/MM_i_2 XI31/XI1/XI44/XI25/Z_NEG XI31/XI1/NET16
+ XI31/XI1/XI44/XI25/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI25/MM_i_3 XI31/XI1/XI44/XI25/NET_0 XI31/XI1/XI44/S_1<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI44/XI25/MM_i_0 XI31/ARITHMETIC_OUT<12> XI31/XI1/XI44/XI25/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI25/MM_i_11 VDD! XI31/XI1/NET16 XI31/XI1/XI44/XI25/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI25/MM_i_8 VDD! XI31/XI1/XI44/S_0<1> XI31/XI1/XI44/XI25/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI25/MM_i_6 XI31/XI1/XI44/XI25/NET_2 XI31/XI1/NET16
+ XI31/XI1/XI44/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI25/MM_i_9 XI31/XI1/XI44/XI25/NET_3 XI31/XI1/XI44/XI25/X1
+ XI31/XI1/XI44/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI25/MM_i_7 VDD! XI31/XI1/XI44/S_1<1> XI31/XI1/XI44/XI25/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI25/MM_i_1 XI31/ARITHMETIC_OUT<12> XI31/XI1/XI44/XI25/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI26/MM_i_10 VSS! XI31/XI1/NET16 XI31/XI1/XI44/XI26/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI26/MM_i_4 XI31/XI1/XI44/XI26/NET_1 XI31/XI1/XI44/S_0<2> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI26/MM_i_5 XI31/XI1/XI44/XI26/Z_NEG XI31/XI1/XI44/XI26/X1
+ XI31/XI1/XI44/XI26/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI26/MM_i_2 XI31/XI1/XI44/XI26/Z_NEG XI31/XI1/NET16
+ XI31/XI1/XI44/XI26/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI26/MM_i_3 XI31/XI1/XI44/XI26/NET_0 XI31/XI1/XI44/S_1<2> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI44/XI26/MM_i_0 XI31/ARITHMETIC_OUT<13> XI31/XI1/XI44/XI26/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI26/MM_i_11 VDD! XI31/XI1/NET16 XI31/XI1/XI44/XI26/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI26/MM_i_8 VDD! XI31/XI1/XI44/S_0<2> XI31/XI1/XI44/XI26/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI26/MM_i_6 XI31/XI1/XI44/XI26/NET_2 XI31/XI1/NET16
+ XI31/XI1/XI44/XI26/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI26/MM_i_9 XI31/XI1/XI44/XI26/NET_3 XI31/XI1/XI44/XI26/X1
+ XI31/XI1/XI44/XI26/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI26/MM_i_7 VDD! XI31/XI1/XI44/S_1<2> XI31/XI1/XI44/XI26/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI26/MM_i_1 XI31/ARITHMETIC_OUT<13> XI31/XI1/XI44/XI26/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI24/MM_i_10 VSS! XI31/XI1/NET16 XI31/XI1/XI44/XI24/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI24/MM_i_4 XI31/XI1/XI44/XI24/NET_1 XI31/XI1/XI44/S_0<3> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI24/MM_i_5 XI31/XI1/XI44/XI24/Z_NEG XI31/XI1/XI44/XI24/X1
+ XI31/XI1/XI44/XI24/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI24/MM_i_2 XI31/XI1/XI44/XI24/Z_NEG XI31/XI1/NET16
+ XI31/XI1/XI44/XI24/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI24/MM_i_3 XI31/XI1/XI44/XI24/NET_0 XI31/XI1/XI44/S_1<3> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI44/XI24/MM_i_0 XI31/ARITHMETIC_OUT<14> XI31/XI1/XI44/XI24/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI24/MM_i_11 VDD! XI31/XI1/NET16 XI31/XI1/XI44/XI24/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI24/MM_i_8 VDD! XI31/XI1/XI44/S_0<3> XI31/XI1/XI44/XI24/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI24/MM_i_6 XI31/XI1/XI44/XI24/NET_2 XI31/XI1/NET16
+ XI31/XI1/XI44/XI24/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI24/MM_i_9 XI31/XI1/XI44/XI24/NET_3 XI31/XI1/XI44/XI24/X1
+ XI31/XI1/XI44/XI24/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI24/MM_i_7 VDD! XI31/XI1/XI44/S_1<3> XI31/XI1/XI44/XI24/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI24/MM_i_1 XI31/ARITHMETIC_OUT<14> XI31/XI1/XI44/XI24/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI35/MM_i_10 VSS! XI31/XI1/NET16 XI31/XI1/XI44/XI35/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI35/MM_i_4 XI31/XI1/XI44/XI35/NET_1 XI31/XI1/XI44/S_0<4> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI35/MM_i_5 XI31/XI1/XI44/XI35/Z_NEG XI31/XI1/XI44/XI35/X1
+ XI31/XI1/XI44/XI35/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI35/MM_i_2 XI31/XI1/XI44/XI35/Z_NEG XI31/XI1/NET16
+ XI31/XI1/XI44/XI35/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI35/MM_i_3 XI31/XI1/XI44/XI35/NET_0 XI31/XI1/XI44/S_1<4> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI44/XI35/MM_i_0 ARITHMETIC_OUT<15> XI31/XI1/XI44/XI35/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI35/MM_i_11 VDD! XI31/XI1/NET16 XI31/XI1/XI44/XI35/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI35/MM_i_8 VDD! XI31/XI1/XI44/S_0<4> XI31/XI1/XI44/XI35/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI35/MM_i_6 XI31/XI1/XI44/XI35/NET_2 XI31/XI1/NET16
+ XI31/XI1/XI44/XI35/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI35/MM_i_9 XI31/XI1/XI44/XI35/NET_3 XI31/XI1/XI44/XI35/X1
+ XI31/XI1/XI44/XI35/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI35/MM_i_7 VDD! XI31/XI1/XI44/S_1<4> XI31/XI1/XI44/XI35/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI35/MM_i_1 ARITHMETIC_OUT<15> XI31/XI1/XI44/XI35/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI18/MM_i_10 VSS! XI31/XI1/NET16 XI31/XI1/XI44/XI18/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI18/MM_i_4 XI31/XI1/XI44/XI18/NET_1 XI31/XI1/XI44/CO_0 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI18/MM_i_5 XI31/XI1/XI44/XI18/Z_NEG XI31/XI1/XI44/XI18/X1
+ XI31/XI1/XI44/XI18/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI18/MM_i_2 XI31/XI1/XI44/XI18/Z_NEG XI31/XI1/NET16
+ XI31/XI1/XI44/XI18/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI18/MM_i_3 XI31/XI1/XI44/XI18/NET_0 XI31/XI1/XI44/CO_1 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI44/XI18/MM_i_0 CO XI31/XI1/XI44/XI18/Z_NEG VSS! VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI18/MM_i_11 VDD! XI31/XI1/NET16 XI31/XI1/XI44/XI18/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI18/MM_i_8 VDD! XI31/XI1/XI44/CO_0 XI31/XI1/XI44/XI18/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI18/MM_i_6 XI31/XI1/XI44/XI18/NET_2 XI31/XI1/NET16
+ XI31/XI1/XI44/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI18/MM_i_9 XI31/XI1/XI44/XI18/NET_3 XI31/XI1/XI44/XI18/X1
+ XI31/XI1/XI44/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI18/MM_i_7 VDD! XI31/XI1/XI44/CO_1 XI31/XI1/XI44/XI18/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI18/MM_i_1 CO XI31/XI1/XI44/XI18/Z_NEG VDD! VDD! PMOS_VTL
+ L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI9/MM_i_0 XI31/XI1/XI44/XI9/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI9/MM_i_7 VSS! OP0<11> XI31/XI1/XI44/XI9/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI44/XI9/MM_i_13 XI31/XI1/XI44/OP0_TEMP<0> XI31/XI1/XI44/XI9/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI44/XI9/MM_i_19 XI31/XI1/XI44/XI9/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI44/OP0_TEMP<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI44/XI9/MM_i_24 VSS! OP0<11> XI31/XI1/XI44/XI9/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI9/MM_i_30 XI31/XI1/XI44/XI9/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI44/XI9/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI9/MM_i_35 VDD! OP0<11> XI31/XI1/XI44/XI9/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI44/XI9/MM_i_41 XI31/XI1/XI44/XI9/NET_003 XI31/XI1/XI44/XI9/NET_000
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI1/XI44/XI9/MM_i_47 XI31/XI1/XI44/OP0_TEMP<0> CTRL_BUFF<0>
+ XI31/XI1/XI44/XI9/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI44/XI9/MM_i_53 XI31/XI1/XI44/XI9/NET_003 OP0<11>
+ XI31/XI1/XI44/OP0_TEMP<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI10/MM_i_0 XI31/XI1/XI44/XI10/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI10/MM_i_7 VSS! OP0<12> XI31/XI1/XI44/XI10/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI44/XI10/MM_i_13 XI31/XI1/XI44/OP0_TEMP<1> XI31/XI1/XI44/XI10/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI44/XI10/MM_i_19 XI31/XI1/XI44/XI10/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI44/OP0_TEMP<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI44/XI10/MM_i_24 VSS! OP0<12> XI31/XI1/XI44/XI10/NET_001 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI10/MM_i_30 XI31/XI1/XI44/XI10/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI44/XI10/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI10/MM_i_35 VDD! OP0<12> XI31/XI1/XI44/XI10/NET_002 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI44/XI10/MM_i_41 XI31/XI1/XI44/XI10/NET_003
+ XI31/XI1/XI44/XI10/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI44/XI10/MM_i_47 XI31/XI1/XI44/OP0_TEMP<1> CTRL_BUFF<0>
+ XI31/XI1/XI44/XI10/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI44/XI10/MM_i_53 XI31/XI1/XI44/XI10/NET_003 OP0<12>
+ XI31/XI1/XI44/OP0_TEMP<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI11/MM_i_0 XI31/XI1/XI44/XI11/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI11/MM_i_7 VSS! OP0<13> XI31/XI1/XI44/XI11/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI44/XI11/MM_i_13 XI31/XI1/XI44/OP0_TEMP<2> XI31/XI1/XI44/XI11/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI44/XI11/MM_i_19 XI31/XI1/XI44/XI11/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI44/OP0_TEMP<2> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI44/XI11/MM_i_24 VSS! OP0<13> XI31/XI1/XI44/XI11/NET_001 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI11/MM_i_30 XI31/XI1/XI44/XI11/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI44/XI11/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI11/MM_i_35 VDD! OP0<13> XI31/XI1/XI44/XI11/NET_002 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI44/XI11/MM_i_41 XI31/XI1/XI44/XI11/NET_003
+ XI31/XI1/XI44/XI11/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI44/XI11/MM_i_47 XI31/XI1/XI44/OP0_TEMP<2> CTRL_BUFF<0>
+ XI31/XI1/XI44/XI11/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI44/XI11/MM_i_53 XI31/XI1/XI44/XI11/NET_003 OP0<13>
+ XI31/XI1/XI44/OP0_TEMP<2> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI12/MM_i_0 XI31/XI1/XI44/XI12/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI12/MM_i_7 VSS! OP0<14> XI31/XI1/XI44/XI12/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI44/XI12/MM_i_13 XI31/XI1/XI44/OP0_TEMP<3> XI31/XI1/XI44/XI12/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI44/XI12/MM_i_19 XI31/XI1/XI44/XI12/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI44/OP0_TEMP<3> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI44/XI12/MM_i_24 VSS! OP0<14> XI31/XI1/XI44/XI12/NET_001 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI12/MM_i_30 XI31/XI1/XI44/XI12/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI44/XI12/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI12/MM_i_35 VDD! OP0<14> XI31/XI1/XI44/XI12/NET_002 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI44/XI12/MM_i_41 XI31/XI1/XI44/XI12/NET_003
+ XI31/XI1/XI44/XI12/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI44/XI12/MM_i_47 XI31/XI1/XI44/OP0_TEMP<3> CTRL_BUFF<0>
+ XI31/XI1/XI44/XI12/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI44/XI12/MM_i_53 XI31/XI1/XI44/XI12/NET_003 OP0<14>
+ XI31/XI1/XI44/OP0_TEMP<3> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI34/MM_i_0 XI31/XI1/XI44/XI34/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI34/MM_i_7 VSS! OP0<15> XI31/XI1/XI44/XI34/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI44/XI34/MM_i_13 OP0_TEMP<15> XI31/XI1/XI44/XI34/NET_000 VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06
mXI31/XI1/XI44/XI34/MM_i_19 XI31/XI1/XI44/XI34/NET_001 CTRL_BUFF<0> OP0_TEMP<15>
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI34/MM_i_24 VSS! OP0<15> XI31/XI1/XI44/XI34/NET_001 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI34/MM_i_30 XI31/XI1/XI44/XI34/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI44/XI34/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI34/MM_i_35 VDD! OP0<15> XI31/XI1/XI44/XI34/NET_002 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI44/XI34/MM_i_41 XI31/XI1/XI44/XI34/NET_003
+ XI31/XI1/XI44/XI34/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI44/XI34/MM_i_47 OP0_TEMP<15> CTRL_BUFF<0> XI31/XI1/XI44/XI34/NET_003
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI34/MM_i_53 XI31/XI1/XI44/XI34/NET_003 OP0<15> OP0_TEMP<15> VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI5/MM_instance_159 XI31/XI1/XI44/NET36 XI31/XI1/XI44/XI5/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI5/MM_instance_166 VSS! OP1<11> XI31/XI1/XI44/XI5/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_170 XI31/XI1/XI44/XI5/NET_000
+ XI31/XI1/XI44/OP0_TEMP<0> XI31/XI1/XI44/XI5/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_176 XI31/XI1/XI44/XI5/NET_001 VDD!
+ XI31/XI1/XI44/XI5/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI5/MM_instance_188 XI31/XI1/XI44/XI5/NET_002
+ XI31/XI1/XI44/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_182 VSS! OP1<11> XI31/XI1/XI44/XI5/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI5/MM_instance_227 XI31/XI1/XI44/XI5/NET_006 OP1<11> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI5/MM_instance_215 VSS! VDD! XI31/XI1/XI44/XI5/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_221 XI31/XI1/XI44/XI5/NET_006
+ XI31/XI1/XI44/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_209 XI31/XI1/XI44/XI5/NET_005
+ XI31/XI1/XI44/XI5/NET_001 XI31/XI1/XI44/XI5/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_203 XI31/XI1/XI44/XI5/NET_004 VDD!
+ XI31/XI1/XI44/XI5/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI5/MM_instance_199 XI31/XI1/XI44/XI5/NET_003 OP1<11>
+ XI31/XI1/XI44/XI5/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<0>
+ XI31/XI1/XI44/XI5/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI5/MM_instance_233 XI31/XI1/XI44/S_1<0>
+ XI31/XI1/XI44/XI5/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI5/MM_instance_239 XI31/XI1/XI44/NET36 XI31/XI1/XI44/XI5/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI5/MM_instance_246 VDD! OP1<11> XI31/XI1/XI44/XI5/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_251 XI31/XI1/XI44/XI5/NET_007
+ XI31/XI1/XI44/OP0_TEMP<0> XI31/XI1/XI44/XI5/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_257 XI31/XI1/XI44/XI5/NET_001 VDD!
+ XI31/XI1/XI44/XI5/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI5/MM_instance_269 XI31/XI1/XI44/XI5/NET_008
+ XI31/XI1/XI44/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_263 VDD! OP1<11> XI31/XI1/XI44/XI5/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI5/MM_instance_309 XI31/XI1/XI44/XI5/NET_011 OP1<11> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI5/MM_instance_297 VDD! VDD! XI31/XI1/XI44/XI5/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_303 XI31/XI1/XI44/XI5/NET_011
+ XI31/XI1/XI44/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_290 XI31/XI1/XI44/XI5/NET_005
+ XI31/XI1/XI44/XI5/NET_001 XI31/XI1/XI44/XI5/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_284 XI31/XI1/XI44/XI5/NET_010 VDD!
+ XI31/XI1/XI44/XI5/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI5/MM_instance_280 XI31/XI1/XI44/XI5/NET_009 OP1<11>
+ XI31/XI1/XI44/XI5/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<0>
+ XI31/XI1/XI44/XI5/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI5/MM_instance_315 XI31/XI1/XI44/S_1<0>
+ XI31/XI1/XI44/XI5/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI0/MM_instance_159 XI31/XI1/XI44/NET16 XI31/XI1/XI44/XI0/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI0/MM_instance_166 VSS! OP1<11> XI31/XI1/XI44/XI0/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_170 XI31/XI1/XI44/XI0/NET_000
+ XI31/XI1/XI44/OP0_TEMP<0> XI31/XI1/XI44/XI0/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_176 XI31/XI1/XI44/XI0/NET_001 VSS!
+ XI31/XI1/XI44/XI0/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI0/MM_instance_188 XI31/XI1/XI44/XI0/NET_002
+ XI31/XI1/XI44/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_182 VSS! OP1<11> XI31/XI1/XI44/XI0/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI0/MM_instance_227 XI31/XI1/XI44/XI0/NET_006 OP1<11> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI0/MM_instance_215 VSS! VSS! XI31/XI1/XI44/XI0/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_221 XI31/XI1/XI44/XI0/NET_006
+ XI31/XI1/XI44/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_209 XI31/XI1/XI44/XI0/NET_005
+ XI31/XI1/XI44/XI0/NET_001 XI31/XI1/XI44/XI0/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_203 XI31/XI1/XI44/XI0/NET_004 VSS!
+ XI31/XI1/XI44/XI0/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI0/MM_instance_199 XI31/XI1/XI44/XI0/NET_003 OP1<11>
+ XI31/XI1/XI44/XI0/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<0>
+ XI31/XI1/XI44/XI0/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI0/MM_instance_233 XI31/XI1/XI44/S_0<0>
+ XI31/XI1/XI44/XI0/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI0/MM_instance_239 XI31/XI1/XI44/NET16 XI31/XI1/XI44/XI0/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI0/MM_instance_246 VDD! OP1<11> XI31/XI1/XI44/XI0/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_251 XI31/XI1/XI44/XI0/NET_007
+ XI31/XI1/XI44/OP0_TEMP<0> XI31/XI1/XI44/XI0/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_257 XI31/XI1/XI44/XI0/NET_001 VSS!
+ XI31/XI1/XI44/XI0/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI0/MM_instance_269 XI31/XI1/XI44/XI0/NET_008
+ XI31/XI1/XI44/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_263 VDD! OP1<11> XI31/XI1/XI44/XI0/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI0/MM_instance_309 XI31/XI1/XI44/XI0/NET_011 OP1<11> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI0/MM_instance_297 VDD! VSS! XI31/XI1/XI44/XI0/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_303 XI31/XI1/XI44/XI0/NET_011
+ XI31/XI1/XI44/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_290 XI31/XI1/XI44/XI0/NET_005
+ XI31/XI1/XI44/XI0/NET_001 XI31/XI1/XI44/XI0/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_284 XI31/XI1/XI44/XI0/NET_010 VSS!
+ XI31/XI1/XI44/XI0/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI0/MM_instance_280 XI31/XI1/XI44/XI0/NET_009 OP1<11>
+ XI31/XI1/XI44/XI0/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<0>
+ XI31/XI1/XI44/XI0/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI0/MM_instance_315 XI31/XI1/XI44/S_0<0>
+ XI31/XI1/XI44/XI0/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI6/MM_instance_159 XI31/XI1/XI44/NET41 XI31/XI1/XI44/XI6/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI6/MM_instance_166 VSS! OP1<12> XI31/XI1/XI44/XI6/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_170 XI31/XI1/XI44/XI6/NET_000
+ XI31/XI1/XI44/OP0_TEMP<1> XI31/XI1/XI44/XI6/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_176 XI31/XI1/XI44/XI6/NET_001 XI31/XI1/XI44/NET36
+ XI31/XI1/XI44/XI6/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI6/MM_instance_188 XI31/XI1/XI44/XI6/NET_002
+ XI31/XI1/XI44/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_182 VSS! OP1<12> XI31/XI1/XI44/XI6/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI6/MM_instance_227 XI31/XI1/XI44/XI6/NET_006 OP1<12> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI6/MM_instance_215 VSS! XI31/XI1/XI44/NET36
+ XI31/XI1/XI44/XI6/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_221 XI31/XI1/XI44/XI6/NET_006
+ XI31/XI1/XI44/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_209 XI31/XI1/XI44/XI6/NET_005
+ XI31/XI1/XI44/XI6/NET_001 XI31/XI1/XI44/XI6/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_203 XI31/XI1/XI44/XI6/NET_004 XI31/XI1/XI44/NET36
+ XI31/XI1/XI44/XI6/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI6/MM_instance_199 XI31/XI1/XI44/XI6/NET_003 OP1<12>
+ XI31/XI1/XI44/XI6/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<1>
+ XI31/XI1/XI44/XI6/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI6/MM_instance_233 XI31/XI1/XI44/S_1<1>
+ XI31/XI1/XI44/XI6/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI6/MM_instance_239 XI31/XI1/XI44/NET41 XI31/XI1/XI44/XI6/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI6/MM_instance_246 VDD! OP1<12> XI31/XI1/XI44/XI6/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_251 XI31/XI1/XI44/XI6/NET_007
+ XI31/XI1/XI44/OP0_TEMP<1> XI31/XI1/XI44/XI6/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_257 XI31/XI1/XI44/XI6/NET_001 XI31/XI1/XI44/NET36
+ XI31/XI1/XI44/XI6/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI6/MM_instance_269 XI31/XI1/XI44/XI6/NET_008
+ XI31/XI1/XI44/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_263 VDD! OP1<12> XI31/XI1/XI44/XI6/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI6/MM_instance_309 XI31/XI1/XI44/XI6/NET_011 OP1<12> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI6/MM_instance_297 VDD! XI31/XI1/XI44/NET36
+ XI31/XI1/XI44/XI6/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_303 XI31/XI1/XI44/XI6/NET_011
+ XI31/XI1/XI44/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_290 XI31/XI1/XI44/XI6/NET_005
+ XI31/XI1/XI44/XI6/NET_001 XI31/XI1/XI44/XI6/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_284 XI31/XI1/XI44/XI6/NET_010 XI31/XI1/XI44/NET36
+ XI31/XI1/XI44/XI6/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI6/MM_instance_280 XI31/XI1/XI44/XI6/NET_009 OP1<12>
+ XI31/XI1/XI44/XI6/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<1>
+ XI31/XI1/XI44/XI6/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI6/MM_instance_315 XI31/XI1/XI44/S_1<1>
+ XI31/XI1/XI44/XI6/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI1/MM_instance_159 XI31/XI1/XI44/NET21 XI31/XI1/XI44/XI1/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI1/MM_instance_166 VSS! OP1<12> XI31/XI1/XI44/XI1/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_170 XI31/XI1/XI44/XI1/NET_000
+ XI31/XI1/XI44/OP0_TEMP<1> XI31/XI1/XI44/XI1/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_176 XI31/XI1/XI44/XI1/NET_001 XI31/XI1/XI44/NET16
+ XI31/XI1/XI44/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI1/MM_instance_188 XI31/XI1/XI44/XI1/NET_002
+ XI31/XI1/XI44/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_182 VSS! OP1<12> XI31/XI1/XI44/XI1/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI1/MM_instance_227 XI31/XI1/XI44/XI1/NET_006 OP1<12> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI1/MM_instance_215 VSS! XI31/XI1/XI44/NET16
+ XI31/XI1/XI44/XI1/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_221 XI31/XI1/XI44/XI1/NET_006
+ XI31/XI1/XI44/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_209 XI31/XI1/XI44/XI1/NET_005
+ XI31/XI1/XI44/XI1/NET_001 XI31/XI1/XI44/XI1/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_203 XI31/XI1/XI44/XI1/NET_004 XI31/XI1/XI44/NET16
+ XI31/XI1/XI44/XI1/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI1/MM_instance_199 XI31/XI1/XI44/XI1/NET_003 OP1<12>
+ XI31/XI1/XI44/XI1/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<1>
+ XI31/XI1/XI44/XI1/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI1/MM_instance_233 XI31/XI1/XI44/S_0<1>
+ XI31/XI1/XI44/XI1/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI1/MM_instance_239 XI31/XI1/XI44/NET21 XI31/XI1/XI44/XI1/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI1/MM_instance_246 VDD! OP1<12> XI31/XI1/XI44/XI1/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_251 XI31/XI1/XI44/XI1/NET_007
+ XI31/XI1/XI44/OP0_TEMP<1> XI31/XI1/XI44/XI1/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_257 XI31/XI1/XI44/XI1/NET_001 XI31/XI1/XI44/NET16
+ XI31/XI1/XI44/XI1/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI1/MM_instance_269 XI31/XI1/XI44/XI1/NET_008
+ XI31/XI1/XI44/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_263 VDD! OP1<12> XI31/XI1/XI44/XI1/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI1/MM_instance_309 XI31/XI1/XI44/XI1/NET_011 OP1<12> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI1/MM_instance_297 VDD! XI31/XI1/XI44/NET16
+ XI31/XI1/XI44/XI1/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_303 XI31/XI1/XI44/XI1/NET_011
+ XI31/XI1/XI44/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_290 XI31/XI1/XI44/XI1/NET_005
+ XI31/XI1/XI44/XI1/NET_001 XI31/XI1/XI44/XI1/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_284 XI31/XI1/XI44/XI1/NET_010 XI31/XI1/XI44/NET16
+ XI31/XI1/XI44/XI1/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI1/MM_instance_280 XI31/XI1/XI44/XI1/NET_009 OP1<12>
+ XI31/XI1/XI44/XI1/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<1>
+ XI31/XI1/XI44/XI1/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI1/MM_instance_315 XI31/XI1/XI44/S_0<1>
+ XI31/XI1/XI44/XI1/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI7/MM_instance_159 XI31/XI1/XI44/NET46 XI31/XI1/XI44/XI7/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI7/MM_instance_166 VSS! OP1<13> XI31/XI1/XI44/XI7/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_170 XI31/XI1/XI44/XI7/NET_000
+ XI31/XI1/XI44/OP0_TEMP<2> XI31/XI1/XI44/XI7/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_176 XI31/XI1/XI44/XI7/NET_001 XI31/XI1/XI44/NET41
+ XI31/XI1/XI44/XI7/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI7/MM_instance_188 XI31/XI1/XI44/XI7/NET_002
+ XI31/XI1/XI44/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_182 VSS! OP1<13> XI31/XI1/XI44/XI7/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI7/MM_instance_227 XI31/XI1/XI44/XI7/NET_006 OP1<13> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI7/MM_instance_215 VSS! XI31/XI1/XI44/NET41
+ XI31/XI1/XI44/XI7/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_221 XI31/XI1/XI44/XI7/NET_006
+ XI31/XI1/XI44/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_209 XI31/XI1/XI44/XI7/NET_005
+ XI31/XI1/XI44/XI7/NET_001 XI31/XI1/XI44/XI7/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_203 XI31/XI1/XI44/XI7/NET_004 XI31/XI1/XI44/NET41
+ XI31/XI1/XI44/XI7/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI7/MM_instance_199 XI31/XI1/XI44/XI7/NET_003 OP1<13>
+ XI31/XI1/XI44/XI7/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<2>
+ XI31/XI1/XI44/XI7/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI7/MM_instance_233 XI31/XI1/XI44/S_1<2>
+ XI31/XI1/XI44/XI7/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI7/MM_instance_239 XI31/XI1/XI44/NET46 XI31/XI1/XI44/XI7/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI7/MM_instance_246 VDD! OP1<13> XI31/XI1/XI44/XI7/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_251 XI31/XI1/XI44/XI7/NET_007
+ XI31/XI1/XI44/OP0_TEMP<2> XI31/XI1/XI44/XI7/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_257 XI31/XI1/XI44/XI7/NET_001 XI31/XI1/XI44/NET41
+ XI31/XI1/XI44/XI7/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI7/MM_instance_269 XI31/XI1/XI44/XI7/NET_008
+ XI31/XI1/XI44/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_263 VDD! OP1<13> XI31/XI1/XI44/XI7/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI7/MM_instance_309 XI31/XI1/XI44/XI7/NET_011 OP1<13> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI7/MM_instance_297 VDD! XI31/XI1/XI44/NET41
+ XI31/XI1/XI44/XI7/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_303 XI31/XI1/XI44/XI7/NET_011
+ XI31/XI1/XI44/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_290 XI31/XI1/XI44/XI7/NET_005
+ XI31/XI1/XI44/XI7/NET_001 XI31/XI1/XI44/XI7/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_284 XI31/XI1/XI44/XI7/NET_010 XI31/XI1/XI44/NET41
+ XI31/XI1/XI44/XI7/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI7/MM_instance_280 XI31/XI1/XI44/XI7/NET_009 OP1<13>
+ XI31/XI1/XI44/XI7/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<2>
+ XI31/XI1/XI44/XI7/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI7/MM_instance_315 XI31/XI1/XI44/S_1<2>
+ XI31/XI1/XI44/XI7/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI2/MM_instance_159 XI31/XI1/XI44/NET26 XI31/XI1/XI44/XI2/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI2/MM_instance_166 VSS! OP1<13> XI31/XI1/XI44/XI2/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_170 XI31/XI1/XI44/XI2/NET_000
+ XI31/XI1/XI44/OP0_TEMP<2> XI31/XI1/XI44/XI2/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_176 XI31/XI1/XI44/XI2/NET_001 XI31/XI1/XI44/NET21
+ XI31/XI1/XI44/XI2/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI2/MM_instance_188 XI31/XI1/XI44/XI2/NET_002
+ XI31/XI1/XI44/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_182 VSS! OP1<13> XI31/XI1/XI44/XI2/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI2/MM_instance_227 XI31/XI1/XI44/XI2/NET_006 OP1<13> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI2/MM_instance_215 VSS! XI31/XI1/XI44/NET21
+ XI31/XI1/XI44/XI2/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_221 XI31/XI1/XI44/XI2/NET_006
+ XI31/XI1/XI44/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_209 XI31/XI1/XI44/XI2/NET_005
+ XI31/XI1/XI44/XI2/NET_001 XI31/XI1/XI44/XI2/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_203 XI31/XI1/XI44/XI2/NET_004 XI31/XI1/XI44/NET21
+ XI31/XI1/XI44/XI2/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI2/MM_instance_199 XI31/XI1/XI44/XI2/NET_003 OP1<13>
+ XI31/XI1/XI44/XI2/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<2>
+ XI31/XI1/XI44/XI2/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI2/MM_instance_233 XI31/XI1/XI44/S_0<2>
+ XI31/XI1/XI44/XI2/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI2/MM_instance_239 XI31/XI1/XI44/NET26 XI31/XI1/XI44/XI2/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI2/MM_instance_246 VDD! OP1<13> XI31/XI1/XI44/XI2/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_251 XI31/XI1/XI44/XI2/NET_007
+ XI31/XI1/XI44/OP0_TEMP<2> XI31/XI1/XI44/XI2/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_257 XI31/XI1/XI44/XI2/NET_001 XI31/XI1/XI44/NET21
+ XI31/XI1/XI44/XI2/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI2/MM_instance_269 XI31/XI1/XI44/XI2/NET_008
+ XI31/XI1/XI44/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_263 VDD! OP1<13> XI31/XI1/XI44/XI2/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI2/MM_instance_309 XI31/XI1/XI44/XI2/NET_011 OP1<13> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI2/MM_instance_297 VDD! XI31/XI1/XI44/NET21
+ XI31/XI1/XI44/XI2/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_303 XI31/XI1/XI44/XI2/NET_011
+ XI31/XI1/XI44/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_290 XI31/XI1/XI44/XI2/NET_005
+ XI31/XI1/XI44/XI2/NET_001 XI31/XI1/XI44/XI2/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_284 XI31/XI1/XI44/XI2/NET_010 XI31/XI1/XI44/NET21
+ XI31/XI1/XI44/XI2/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI2/MM_instance_280 XI31/XI1/XI44/XI2/NET_009 OP1<13>
+ XI31/XI1/XI44/XI2/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<2>
+ XI31/XI1/XI44/XI2/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI2/MM_instance_315 XI31/XI1/XI44/S_0<2>
+ XI31/XI1/XI44/XI2/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI8/MM_instance_159 XI31/XI1/XI44/NET1 XI31/XI1/XI44/XI8/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI8/MM_instance_166 VSS! OP1<14> XI31/XI1/XI44/XI8/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_170 XI31/XI1/XI44/XI8/NET_000
+ XI31/XI1/XI44/OP0_TEMP<3> XI31/XI1/XI44/XI8/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_176 XI31/XI1/XI44/XI8/NET_001 XI31/XI1/XI44/NET46
+ XI31/XI1/XI44/XI8/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI8/MM_instance_188 XI31/XI1/XI44/XI8/NET_002
+ XI31/XI1/XI44/OP0_TEMP<3> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_182 VSS! OP1<14> XI31/XI1/XI44/XI8/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI8/MM_instance_227 XI31/XI1/XI44/XI8/NET_006 OP1<14> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI8/MM_instance_215 VSS! XI31/XI1/XI44/NET46
+ XI31/XI1/XI44/XI8/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_221 XI31/XI1/XI44/XI8/NET_006
+ XI31/XI1/XI44/OP0_TEMP<3> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_209 XI31/XI1/XI44/XI8/NET_005
+ XI31/XI1/XI44/XI8/NET_001 XI31/XI1/XI44/XI8/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_203 XI31/XI1/XI44/XI8/NET_004 XI31/XI1/XI44/NET46
+ XI31/XI1/XI44/XI8/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI8/MM_instance_199 XI31/XI1/XI44/XI8/NET_003 OP1<14>
+ XI31/XI1/XI44/XI8/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<3>
+ XI31/XI1/XI44/XI8/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI8/MM_instance_233 XI31/XI1/XI44/S_1<3>
+ XI31/XI1/XI44/XI8/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI8/MM_instance_239 XI31/XI1/XI44/NET1 XI31/XI1/XI44/XI8/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI8/MM_instance_246 VDD! OP1<14> XI31/XI1/XI44/XI8/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_251 XI31/XI1/XI44/XI8/NET_007
+ XI31/XI1/XI44/OP0_TEMP<3> XI31/XI1/XI44/XI8/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_257 XI31/XI1/XI44/XI8/NET_001 XI31/XI1/XI44/NET46
+ XI31/XI1/XI44/XI8/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI8/MM_instance_269 XI31/XI1/XI44/XI8/NET_008
+ XI31/XI1/XI44/OP0_TEMP<3> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_263 VDD! OP1<14> XI31/XI1/XI44/XI8/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI8/MM_instance_309 XI31/XI1/XI44/XI8/NET_011 OP1<14> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI8/MM_instance_297 VDD! XI31/XI1/XI44/NET46
+ XI31/XI1/XI44/XI8/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_303 XI31/XI1/XI44/XI8/NET_011
+ XI31/XI1/XI44/OP0_TEMP<3> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_290 XI31/XI1/XI44/XI8/NET_005
+ XI31/XI1/XI44/XI8/NET_001 XI31/XI1/XI44/XI8/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_284 XI31/XI1/XI44/XI8/NET_010 XI31/XI1/XI44/NET46
+ XI31/XI1/XI44/XI8/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI8/MM_instance_280 XI31/XI1/XI44/XI8/NET_009 OP1<14>
+ XI31/XI1/XI44/XI8/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<3>
+ XI31/XI1/XI44/XI8/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI8/MM_instance_315 XI31/XI1/XI44/S_1<3>
+ XI31/XI1/XI44/XI8/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI3/MM_instance_159 XI31/XI1/XI44/NET2 XI31/XI1/XI44/XI3/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI44/XI3/MM_instance_166 VSS! OP1<14> XI31/XI1/XI44/XI3/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_170 XI31/XI1/XI44/XI3/NET_000
+ XI31/XI1/XI44/OP0_TEMP<3> XI31/XI1/XI44/XI3/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_176 XI31/XI1/XI44/XI3/NET_001 XI31/XI1/XI44/NET26
+ XI31/XI1/XI44/XI3/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI3/MM_instance_188 XI31/XI1/XI44/XI3/NET_002
+ XI31/XI1/XI44/OP0_TEMP<3> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_182 VSS! OP1<14> XI31/XI1/XI44/XI3/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI3/MM_instance_227 XI31/XI1/XI44/XI3/NET_006 OP1<14> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI3/MM_instance_215 VSS! XI31/XI1/XI44/NET26
+ XI31/XI1/XI44/XI3/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_221 XI31/XI1/XI44/XI3/NET_006
+ XI31/XI1/XI44/OP0_TEMP<3> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_209 XI31/XI1/XI44/XI3/NET_005
+ XI31/XI1/XI44/XI3/NET_001 XI31/XI1/XI44/XI3/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_203 XI31/XI1/XI44/XI3/NET_004 XI31/XI1/XI44/NET26
+ XI31/XI1/XI44/XI3/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI3/MM_instance_199 XI31/XI1/XI44/XI3/NET_003 OP1<14>
+ XI31/XI1/XI44/XI3/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_194 VSS! XI31/XI1/XI44/OP0_TEMP<3>
+ XI31/XI1/XI44/XI3/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI3/MM_instance_233 XI31/XI1/XI44/S_0<3>
+ XI31/XI1/XI44/XI3/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI3/MM_instance_239 XI31/XI1/XI44/NET2 XI31/XI1/XI44/XI3/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI44/XI3/MM_instance_246 VDD! OP1<14> XI31/XI1/XI44/XI3/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_251 XI31/XI1/XI44/XI3/NET_007
+ XI31/XI1/XI44/OP0_TEMP<3> XI31/XI1/XI44/XI3/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_257 XI31/XI1/XI44/XI3/NET_001 XI31/XI1/XI44/NET26
+ XI31/XI1/XI44/XI3/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI3/MM_instance_269 XI31/XI1/XI44/XI3/NET_008
+ XI31/XI1/XI44/OP0_TEMP<3> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_263 VDD! OP1<14> XI31/XI1/XI44/XI3/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI3/MM_instance_309 XI31/XI1/XI44/XI3/NET_011 OP1<14> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI3/MM_instance_297 VDD! XI31/XI1/XI44/NET26
+ XI31/XI1/XI44/XI3/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_303 XI31/XI1/XI44/XI3/NET_011
+ XI31/XI1/XI44/OP0_TEMP<3> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_290 XI31/XI1/XI44/XI3/NET_005
+ XI31/XI1/XI44/XI3/NET_001 XI31/XI1/XI44/XI3/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_284 XI31/XI1/XI44/XI3/NET_010 XI31/XI1/XI44/NET26
+ XI31/XI1/XI44/XI3/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI3/MM_instance_280 XI31/XI1/XI44/XI3/NET_009 OP1<14>
+ XI31/XI1/XI44/XI3/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_275 VDD! XI31/XI1/XI44/OP0_TEMP<3>
+ XI31/XI1/XI44/XI3/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI3/MM_instance_315 XI31/XI1/XI44/S_0<3>
+ XI31/XI1/XI44/XI3/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI32/MM_instance_159 XI31/XI1/XI44/CO_1
+ XI31/XI1/XI44/XI32/NET_001 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI32/MM_instance_166 VSS! OP1<15> XI31/XI1/XI44/XI32/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_170 XI31/XI1/XI44/XI32/NET_000 OP0_TEMP<15>
+ XI31/XI1/XI44/XI32/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_176 XI31/XI1/XI44/XI32/NET_001
+ XI31/XI1/XI44/NET1 XI31/XI1/XI44/XI32/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI32/MM_instance_188 XI31/XI1/XI44/XI32/NET_002 OP0_TEMP<15> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_182 VSS! OP1<15> XI31/XI1/XI44/XI32/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI32/MM_instance_227 XI31/XI1/XI44/XI32/NET_006 OP1<15> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI32/MM_instance_215 VSS! XI31/XI1/XI44/NET1
+ XI31/XI1/XI44/XI32/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_221 XI31/XI1/XI44/XI32/NET_006 OP0_TEMP<15> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_209 XI31/XI1/XI44/XI32/NET_005
+ XI31/XI1/XI44/XI32/NET_001 XI31/XI1/XI44/XI32/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_203 XI31/XI1/XI44/XI32/NET_004
+ XI31/XI1/XI44/NET1 XI31/XI1/XI44/XI32/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI32/MM_instance_199 XI31/XI1/XI44/XI32/NET_003 OP1<15>
+ XI31/XI1/XI44/XI32/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_194 VSS! OP0_TEMP<15> XI31/XI1/XI44/XI32/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI32/MM_instance_233 XI31/XI1/XI44/S_1<4>
+ XI31/XI1/XI44/XI32/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI32/MM_instance_239 XI31/XI1/XI44/CO_1
+ XI31/XI1/XI44/XI32/NET_001 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI32/MM_instance_246 VDD! OP1<15> XI31/XI1/XI44/XI32/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_251 XI31/XI1/XI44/XI32/NET_007 OP0_TEMP<15>
+ XI31/XI1/XI44/XI32/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_257 XI31/XI1/XI44/XI32/NET_001
+ XI31/XI1/XI44/NET1 XI31/XI1/XI44/XI32/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI32/MM_instance_269 XI31/XI1/XI44/XI32/NET_008 OP0_TEMP<15> VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_263 VDD! OP1<15> XI31/XI1/XI44/XI32/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI32/MM_instance_309 XI31/XI1/XI44/XI32/NET_011 OP1<15> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI32/MM_instance_297 VDD! XI31/XI1/XI44/NET1
+ XI31/XI1/XI44/XI32/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_303 XI31/XI1/XI44/XI32/NET_011 OP0_TEMP<15> VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_290 XI31/XI1/XI44/XI32/NET_005
+ XI31/XI1/XI44/XI32/NET_001 XI31/XI1/XI44/XI32/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_284 XI31/XI1/XI44/XI32/NET_010
+ XI31/XI1/XI44/NET1 XI31/XI1/XI44/XI32/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI32/MM_instance_280 XI31/XI1/XI44/XI32/NET_009 OP1<15>
+ XI31/XI1/XI44/XI32/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_275 VDD! OP0_TEMP<15> XI31/XI1/XI44/XI32/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI32/MM_instance_315 XI31/XI1/XI44/S_1<4>
+ XI31/XI1/XI44/XI32/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI33/MM_instance_159 XI31/XI1/XI44/CO_0
+ XI31/XI1/XI44/XI33/NET_001 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI33/MM_instance_166 VSS! OP1<15> XI31/XI1/XI44/XI33/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_170 XI31/XI1/XI44/XI33/NET_000 OP0_TEMP<15>
+ XI31/XI1/XI44/XI33/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_176 XI31/XI1/XI44/XI33/NET_001
+ XI31/XI1/XI44/NET2 XI31/XI1/XI44/XI33/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI44/XI33/MM_instance_188 XI31/XI1/XI44/XI33/NET_002 OP0_TEMP<15> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_182 VSS! OP1<15> XI31/XI1/XI44/XI33/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI33/MM_instance_227 XI31/XI1/XI44/XI33/NET_006 OP1<15> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI44/XI33/MM_instance_215 VSS! XI31/XI1/XI44/NET2
+ XI31/XI1/XI44/XI33/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_221 XI31/XI1/XI44/XI33/NET_006 OP0_TEMP<15> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_209 XI31/XI1/XI44/XI33/NET_005
+ XI31/XI1/XI44/XI33/NET_001 XI31/XI1/XI44/XI33/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_203 XI31/XI1/XI44/XI33/NET_004
+ XI31/XI1/XI44/NET2 XI31/XI1/XI44/XI33/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07
+ AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI44/XI33/MM_instance_199 XI31/XI1/XI44/XI33/NET_003 OP1<15>
+ XI31/XI1/XI44/XI33/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_194 VSS! OP0_TEMP<15> XI31/XI1/XI44/XI33/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI44/XI33/MM_instance_233 XI31/XI1/XI44/S_0<4>
+ XI31/XI1/XI44/XI33/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI44/XI33/MM_instance_239 XI31/XI1/XI44/CO_0
+ XI31/XI1/XI44/XI33/NET_001 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI44/XI33/MM_instance_246 VDD! OP1<15> XI31/XI1/XI44/XI33/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_251 XI31/XI1/XI44/XI33/NET_007 OP0_TEMP<15>
+ XI31/XI1/XI44/XI33/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_257 XI31/XI1/XI44/XI33/NET_001
+ XI31/XI1/XI44/NET2 XI31/XI1/XI44/XI33/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI44/XI33/MM_instance_269 XI31/XI1/XI44/XI33/NET_008 OP0_TEMP<15> VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_263 VDD! OP1<15> XI31/XI1/XI44/XI33/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI33/MM_instance_309 XI31/XI1/XI44/XI33/NET_011 OP1<15> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI44/XI33/MM_instance_297 VDD! XI31/XI1/XI44/NET2
+ XI31/XI1/XI44/XI33/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_303 XI31/XI1/XI44/XI33/NET_011 OP0_TEMP<15> VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_290 XI31/XI1/XI44/XI33/NET_005
+ XI31/XI1/XI44/XI33/NET_001 XI31/XI1/XI44/XI33/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_284 XI31/XI1/XI44/XI33/NET_010
+ XI31/XI1/XI44/NET2 XI31/XI1/XI44/XI33/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07
+ AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI44/XI33/MM_instance_280 XI31/XI1/XI44/XI33/NET_009 OP1<15>
+ XI31/XI1/XI44/XI33/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_275 VDD! OP0_TEMP<15> XI31/XI1/XI44/XI33/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI44/XI33/MM_instance_315 XI31/XI1/XI44/S_0<4>
+ XI31/XI1/XI44/XI33/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI17/MM_i_10 VSS! XI31/XI1/NET12 XI31/XI1/XI43/XI17/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI17/MM_i_4 XI31/XI1/XI43/XI17/NET_1 XI31/XI1/XI43/S_0<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI17/MM_i_5 XI31/XI1/XI43/XI17/Z_NEG XI31/XI1/XI43/XI17/X1
+ XI31/XI1/XI43/XI17/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI17/MM_i_2 XI31/XI1/XI43/XI17/Z_NEG XI31/XI1/NET12
+ XI31/XI1/XI43/XI17/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI17/MM_i_3 XI31/XI1/XI43/XI17/NET_0 XI31/XI1/XI43/S_1<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI43/XI17/MM_i_0 XI31/ARITHMETIC_OUT<7> XI31/XI1/XI43/XI17/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI17/MM_i_11 VDD! XI31/XI1/NET12 XI31/XI1/XI43/XI17/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI17/MM_i_8 VDD! XI31/XI1/XI43/S_0<0> XI31/XI1/XI43/XI17/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI17/MM_i_6 XI31/XI1/XI43/XI17/NET_2 XI31/XI1/NET12
+ XI31/XI1/XI43/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI17/MM_i_9 XI31/XI1/XI43/XI17/NET_3 XI31/XI1/XI43/XI17/X1
+ XI31/XI1/XI43/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI17/MM_i_7 VDD! XI31/XI1/XI43/S_1<0> XI31/XI1/XI43/XI17/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI17/MM_i_1 XI31/ARITHMETIC_OUT<7> XI31/XI1/XI43/XI17/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI25/MM_i_10 VSS! XI31/XI1/NET12 XI31/XI1/XI43/XI25/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI25/MM_i_4 XI31/XI1/XI43/XI25/NET_1 XI31/XI1/XI43/S_0<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI25/MM_i_5 XI31/XI1/XI43/XI25/Z_NEG XI31/XI1/XI43/XI25/X1
+ XI31/XI1/XI43/XI25/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI25/MM_i_2 XI31/XI1/XI43/XI25/Z_NEG XI31/XI1/NET12
+ XI31/XI1/XI43/XI25/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI25/MM_i_3 XI31/XI1/XI43/XI25/NET_0 XI31/XI1/XI43/S_1<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI43/XI25/MM_i_0 XI31/ARITHMETIC_OUT<8> XI31/XI1/XI43/XI25/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI25/MM_i_11 VDD! XI31/XI1/NET12 XI31/XI1/XI43/XI25/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI25/MM_i_8 VDD! XI31/XI1/XI43/S_0<1> XI31/XI1/XI43/XI25/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI25/MM_i_6 XI31/XI1/XI43/XI25/NET_2 XI31/XI1/NET12
+ XI31/XI1/XI43/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI25/MM_i_9 XI31/XI1/XI43/XI25/NET_3 XI31/XI1/XI43/XI25/X1
+ XI31/XI1/XI43/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI25/MM_i_7 VDD! XI31/XI1/XI43/S_1<1> XI31/XI1/XI43/XI25/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI25/MM_i_1 XI31/ARITHMETIC_OUT<8> XI31/XI1/XI43/XI25/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI26/MM_i_10 VSS! XI31/XI1/NET12 XI31/XI1/XI43/XI26/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI26/MM_i_4 XI31/XI1/XI43/XI26/NET_1 XI31/XI1/XI43/S_0<2> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI26/MM_i_5 XI31/XI1/XI43/XI26/Z_NEG XI31/XI1/XI43/XI26/X1
+ XI31/XI1/XI43/XI26/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI26/MM_i_2 XI31/XI1/XI43/XI26/Z_NEG XI31/XI1/NET12
+ XI31/XI1/XI43/XI26/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI26/MM_i_3 XI31/XI1/XI43/XI26/NET_0 XI31/XI1/XI43/S_1<2> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI43/XI26/MM_i_0 XI31/ARITHMETIC_OUT<9> XI31/XI1/XI43/XI26/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI26/MM_i_11 VDD! XI31/XI1/NET12 XI31/XI1/XI43/XI26/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI26/MM_i_8 VDD! XI31/XI1/XI43/S_0<2> XI31/XI1/XI43/XI26/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI26/MM_i_6 XI31/XI1/XI43/XI26/NET_2 XI31/XI1/NET12
+ XI31/XI1/XI43/XI26/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI26/MM_i_9 XI31/XI1/XI43/XI26/NET_3 XI31/XI1/XI43/XI26/X1
+ XI31/XI1/XI43/XI26/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI26/MM_i_7 VDD! XI31/XI1/XI43/S_1<2> XI31/XI1/XI43/XI26/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI26/MM_i_1 XI31/ARITHMETIC_OUT<9> XI31/XI1/XI43/XI26/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI24/MM_i_10 VSS! XI31/XI1/NET12 XI31/XI1/XI43/XI24/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI24/MM_i_4 XI31/XI1/XI43/XI24/NET_1 XI31/XI1/XI43/S_0<3> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI24/MM_i_5 XI31/XI1/XI43/XI24/Z_NEG XI31/XI1/XI43/XI24/X1
+ XI31/XI1/XI43/XI24/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI24/MM_i_2 XI31/XI1/XI43/XI24/Z_NEG XI31/XI1/NET12
+ XI31/XI1/XI43/XI24/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI24/MM_i_3 XI31/XI1/XI43/XI24/NET_0 XI31/XI1/XI43/S_1<3> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI43/XI24/MM_i_0 XI31/ARITHMETIC_OUT<10> XI31/XI1/XI43/XI24/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI24/MM_i_11 VDD! XI31/XI1/NET12 XI31/XI1/XI43/XI24/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI24/MM_i_8 VDD! XI31/XI1/XI43/S_0<3> XI31/XI1/XI43/XI24/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI24/MM_i_6 XI31/XI1/XI43/XI24/NET_2 XI31/XI1/NET12
+ XI31/XI1/XI43/XI24/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI24/MM_i_9 XI31/XI1/XI43/XI24/NET_3 XI31/XI1/XI43/XI24/X1
+ XI31/XI1/XI43/XI24/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI24/MM_i_7 VDD! XI31/XI1/XI43/S_1<3> XI31/XI1/XI43/XI24/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI24/MM_i_1 XI31/ARITHMETIC_OUT<10> XI31/XI1/XI43/XI24/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI18/MM_i_10 VSS! XI31/XI1/NET12 XI31/XI1/XI43/XI18/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI18/MM_i_4 XI31/XI1/XI43/XI18/NET_1 XI31/XI1/XI43/CO_0 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI18/MM_i_5 XI31/XI1/XI43/XI18/Z_NEG XI31/XI1/XI43/XI18/X1
+ XI31/XI1/XI43/XI18/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI18/MM_i_2 XI31/XI1/XI43/XI18/Z_NEG XI31/XI1/NET12
+ XI31/XI1/XI43/XI18/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI18/MM_i_3 XI31/XI1/XI43/XI18/NET_0 XI31/XI1/XI43/CO_1 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI43/XI18/MM_i_0 XI31/XI1/NET16 XI31/XI1/XI43/XI18/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI18/MM_i_11 VDD! XI31/XI1/NET12 XI31/XI1/XI43/XI18/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI18/MM_i_8 VDD! XI31/XI1/XI43/CO_0 XI31/XI1/XI43/XI18/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI18/MM_i_6 XI31/XI1/XI43/XI18/NET_2 XI31/XI1/NET12
+ XI31/XI1/XI43/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI18/MM_i_9 XI31/XI1/XI43/XI18/NET_3 XI31/XI1/XI43/XI18/X1
+ XI31/XI1/XI43/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI18/MM_i_7 VDD! XI31/XI1/XI43/CO_1 XI31/XI1/XI43/XI18/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI18/MM_i_1 XI31/XI1/NET16 XI31/XI1/XI43/XI18/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI9/MM_i_0 XI31/XI1/XI43/XI9/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI9/MM_i_7 VSS! OP0<7> XI31/XI1/XI43/XI9/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI43/XI9/MM_i_13 XI31/XI1/XI43/OP0_TEMP<0> XI31/XI1/XI43/XI9/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI43/XI9/MM_i_19 XI31/XI1/XI43/XI9/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI43/OP0_TEMP<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI43/XI9/MM_i_24 VSS! OP0<7> XI31/XI1/XI43/XI9/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI9/MM_i_30 XI31/XI1/XI43/XI9/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI43/XI9/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI9/MM_i_35 VDD! OP0<7> XI31/XI1/XI43/XI9/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI43/XI9/MM_i_41 XI31/XI1/XI43/XI9/NET_003 XI31/XI1/XI43/XI9/NET_000
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI1/XI43/XI9/MM_i_47 XI31/XI1/XI43/OP0_TEMP<0> CTRL_BUFF<0>
+ XI31/XI1/XI43/XI9/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI43/XI9/MM_i_53 XI31/XI1/XI43/XI9/NET_003 OP0<7>
+ XI31/XI1/XI43/OP0_TEMP<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI10/MM_i_0 XI31/XI1/XI43/XI10/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI10/MM_i_7 VSS! OP0<8> XI31/XI1/XI43/XI10/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI43/XI10/MM_i_13 XI31/XI1/XI43/OP0_TEMP<1> XI31/XI1/XI43/XI10/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI43/XI10/MM_i_19 XI31/XI1/XI43/XI10/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI43/OP0_TEMP<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI43/XI10/MM_i_24 VSS! OP0<8> XI31/XI1/XI43/XI10/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI10/MM_i_30 XI31/XI1/XI43/XI10/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI43/XI10/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI10/MM_i_35 VDD! OP0<8> XI31/XI1/XI43/XI10/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI43/XI10/MM_i_41 XI31/XI1/XI43/XI10/NET_003
+ XI31/XI1/XI43/XI10/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI43/XI10/MM_i_47 XI31/XI1/XI43/OP0_TEMP<1> CTRL_BUFF<0>
+ XI31/XI1/XI43/XI10/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI43/XI10/MM_i_53 XI31/XI1/XI43/XI10/NET_003 OP0<8>
+ XI31/XI1/XI43/OP0_TEMP<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI11/MM_i_0 XI31/XI1/XI43/XI11/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI11/MM_i_7 VSS! OP0<9> XI31/XI1/XI43/XI11/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI43/XI11/MM_i_13 XI31/XI1/XI43/OP0_TEMP<2> XI31/XI1/XI43/XI11/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI43/XI11/MM_i_19 XI31/XI1/XI43/XI11/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI43/OP0_TEMP<2> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI43/XI11/MM_i_24 VSS! OP0<9> XI31/XI1/XI43/XI11/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI11/MM_i_30 XI31/XI1/XI43/XI11/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI43/XI11/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI11/MM_i_35 VDD! OP0<9> XI31/XI1/XI43/XI11/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI43/XI11/MM_i_41 XI31/XI1/XI43/XI11/NET_003
+ XI31/XI1/XI43/XI11/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI43/XI11/MM_i_47 XI31/XI1/XI43/OP0_TEMP<2> CTRL_BUFF<0>
+ XI31/XI1/XI43/XI11/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI43/XI11/MM_i_53 XI31/XI1/XI43/XI11/NET_003 OP0<9>
+ XI31/XI1/XI43/OP0_TEMP<2> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI12/MM_i_0 XI31/XI1/XI43/XI12/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI12/MM_i_7 VSS! OP0<10> XI31/XI1/XI43/XI12/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI43/XI12/MM_i_13 XI31/XI1/NET18 XI31/XI1/XI43/XI12/NET_000 VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06
mXI31/XI1/XI43/XI12/MM_i_19 XI31/XI1/XI43/XI12/NET_001 CTRL_BUFF<0>
+ XI31/XI1/NET18 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14
+ PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI43/XI12/MM_i_24 VSS! OP0<10> XI31/XI1/XI43/XI12/NET_001 VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI12/MM_i_30 XI31/XI1/XI43/XI12/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI43/XI12/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI12/MM_i_35 VDD! OP0<10> XI31/XI1/XI43/XI12/NET_002 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI43/XI12/MM_i_41 XI31/XI1/XI43/XI12/NET_003
+ XI31/XI1/XI43/XI12/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI43/XI12/MM_i_47 XI31/XI1/NET18 CTRL_BUFF<0>
+ XI31/XI1/XI43/XI12/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI43/XI12/MM_i_53 XI31/XI1/XI43/XI12/NET_003 OP0<10> XI31/XI1/NET18
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI5/MM_instance_159 XI31/XI1/XI43/NET36 XI31/XI1/XI43/XI5/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI5/MM_instance_166 VSS! OP1<7> XI31/XI1/XI43/XI5/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_170 XI31/XI1/XI43/XI5/NET_000
+ XI31/XI1/XI43/OP0_TEMP<0> XI31/XI1/XI43/XI5/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_176 XI31/XI1/XI43/XI5/NET_001 VDD!
+ XI31/XI1/XI43/XI5/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI5/MM_instance_188 XI31/XI1/XI43/XI5/NET_002
+ XI31/XI1/XI43/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_182 VSS! OP1<7> XI31/XI1/XI43/XI5/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI5/MM_instance_227 XI31/XI1/XI43/XI5/NET_006 OP1<7> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI5/MM_instance_215 VSS! VDD! XI31/XI1/XI43/XI5/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_221 XI31/XI1/XI43/XI5/NET_006
+ XI31/XI1/XI43/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_209 XI31/XI1/XI43/XI5/NET_005
+ XI31/XI1/XI43/XI5/NET_001 XI31/XI1/XI43/XI5/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_203 XI31/XI1/XI43/XI5/NET_004 VDD!
+ XI31/XI1/XI43/XI5/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI5/MM_instance_199 XI31/XI1/XI43/XI5/NET_003 OP1<7>
+ XI31/XI1/XI43/XI5/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_194 VSS! XI31/XI1/XI43/OP0_TEMP<0>
+ XI31/XI1/XI43/XI5/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI5/MM_instance_233 XI31/XI1/XI43/S_1<0>
+ XI31/XI1/XI43/XI5/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI5/MM_instance_239 XI31/XI1/XI43/NET36 XI31/XI1/XI43/XI5/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI5/MM_instance_246 VDD! OP1<7> XI31/XI1/XI43/XI5/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_251 XI31/XI1/XI43/XI5/NET_007
+ XI31/XI1/XI43/OP0_TEMP<0> XI31/XI1/XI43/XI5/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_257 XI31/XI1/XI43/XI5/NET_001 VDD!
+ XI31/XI1/XI43/XI5/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI5/MM_instance_269 XI31/XI1/XI43/XI5/NET_008
+ XI31/XI1/XI43/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_263 VDD! OP1<7> XI31/XI1/XI43/XI5/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI5/MM_instance_309 XI31/XI1/XI43/XI5/NET_011 OP1<7> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI5/MM_instance_297 VDD! VDD! XI31/XI1/XI43/XI5/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_303 XI31/XI1/XI43/XI5/NET_011
+ XI31/XI1/XI43/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_290 XI31/XI1/XI43/XI5/NET_005
+ XI31/XI1/XI43/XI5/NET_001 XI31/XI1/XI43/XI5/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_284 XI31/XI1/XI43/XI5/NET_010 VDD!
+ XI31/XI1/XI43/XI5/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI5/MM_instance_280 XI31/XI1/XI43/XI5/NET_009 OP1<7>
+ XI31/XI1/XI43/XI5/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_275 VDD! XI31/XI1/XI43/OP0_TEMP<0>
+ XI31/XI1/XI43/XI5/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI5/MM_instance_315 XI31/XI1/XI43/S_1<0>
+ XI31/XI1/XI43/XI5/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI0/MM_instance_159 XI31/XI1/XI43/NET16 XI31/XI1/XI43/XI0/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI0/MM_instance_166 VSS! OP1<7> XI31/XI1/XI43/XI0/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_170 XI31/XI1/XI43/XI0/NET_000
+ XI31/XI1/XI43/OP0_TEMP<0> XI31/XI1/XI43/XI0/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_176 XI31/XI1/XI43/XI0/NET_001 VSS!
+ XI31/XI1/XI43/XI0/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI0/MM_instance_188 XI31/XI1/XI43/XI0/NET_002
+ XI31/XI1/XI43/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_182 VSS! OP1<7> XI31/XI1/XI43/XI0/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI0/MM_instance_227 XI31/XI1/XI43/XI0/NET_006 OP1<7> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI0/MM_instance_215 VSS! VSS! XI31/XI1/XI43/XI0/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_221 XI31/XI1/XI43/XI0/NET_006
+ XI31/XI1/XI43/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_209 XI31/XI1/XI43/XI0/NET_005
+ XI31/XI1/XI43/XI0/NET_001 XI31/XI1/XI43/XI0/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_203 XI31/XI1/XI43/XI0/NET_004 VSS!
+ XI31/XI1/XI43/XI0/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI0/MM_instance_199 XI31/XI1/XI43/XI0/NET_003 OP1<7>
+ XI31/XI1/XI43/XI0/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_194 VSS! XI31/XI1/XI43/OP0_TEMP<0>
+ XI31/XI1/XI43/XI0/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI0/MM_instance_233 XI31/XI1/XI43/S_0<0>
+ XI31/XI1/XI43/XI0/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI0/MM_instance_239 XI31/XI1/XI43/NET16 XI31/XI1/XI43/XI0/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI0/MM_instance_246 VDD! OP1<7> XI31/XI1/XI43/XI0/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_251 XI31/XI1/XI43/XI0/NET_007
+ XI31/XI1/XI43/OP0_TEMP<0> XI31/XI1/XI43/XI0/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_257 XI31/XI1/XI43/XI0/NET_001 VSS!
+ XI31/XI1/XI43/XI0/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI0/MM_instance_269 XI31/XI1/XI43/XI0/NET_008
+ XI31/XI1/XI43/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_263 VDD! OP1<7> XI31/XI1/XI43/XI0/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI0/MM_instance_309 XI31/XI1/XI43/XI0/NET_011 OP1<7> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI0/MM_instance_297 VDD! VSS! XI31/XI1/XI43/XI0/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_303 XI31/XI1/XI43/XI0/NET_011
+ XI31/XI1/XI43/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_290 XI31/XI1/XI43/XI0/NET_005
+ XI31/XI1/XI43/XI0/NET_001 XI31/XI1/XI43/XI0/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_284 XI31/XI1/XI43/XI0/NET_010 VSS!
+ XI31/XI1/XI43/XI0/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI0/MM_instance_280 XI31/XI1/XI43/XI0/NET_009 OP1<7>
+ XI31/XI1/XI43/XI0/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_275 VDD! XI31/XI1/XI43/OP0_TEMP<0>
+ XI31/XI1/XI43/XI0/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI0/MM_instance_315 XI31/XI1/XI43/S_0<0>
+ XI31/XI1/XI43/XI0/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI6/MM_instance_159 XI31/XI1/XI43/NET41 XI31/XI1/XI43/XI6/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI6/MM_instance_166 VSS! OP1<8> XI31/XI1/XI43/XI6/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_170 XI31/XI1/XI43/XI6/NET_000
+ XI31/XI1/XI43/OP0_TEMP<1> XI31/XI1/XI43/XI6/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_176 XI31/XI1/XI43/XI6/NET_001 XI31/XI1/XI43/NET36
+ XI31/XI1/XI43/XI6/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI6/MM_instance_188 XI31/XI1/XI43/XI6/NET_002
+ XI31/XI1/XI43/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_182 VSS! OP1<8> XI31/XI1/XI43/XI6/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI6/MM_instance_227 XI31/XI1/XI43/XI6/NET_006 OP1<8> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI6/MM_instance_215 VSS! XI31/XI1/XI43/NET36
+ XI31/XI1/XI43/XI6/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_221 XI31/XI1/XI43/XI6/NET_006
+ XI31/XI1/XI43/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_209 XI31/XI1/XI43/XI6/NET_005
+ XI31/XI1/XI43/XI6/NET_001 XI31/XI1/XI43/XI6/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_203 XI31/XI1/XI43/XI6/NET_004 XI31/XI1/XI43/NET36
+ XI31/XI1/XI43/XI6/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI6/MM_instance_199 XI31/XI1/XI43/XI6/NET_003 OP1<8>
+ XI31/XI1/XI43/XI6/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_194 VSS! XI31/XI1/XI43/OP0_TEMP<1>
+ XI31/XI1/XI43/XI6/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI6/MM_instance_233 XI31/XI1/XI43/S_1<1>
+ XI31/XI1/XI43/XI6/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI6/MM_instance_239 XI31/XI1/XI43/NET41 XI31/XI1/XI43/XI6/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI6/MM_instance_246 VDD! OP1<8> XI31/XI1/XI43/XI6/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_251 XI31/XI1/XI43/XI6/NET_007
+ XI31/XI1/XI43/OP0_TEMP<1> XI31/XI1/XI43/XI6/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_257 XI31/XI1/XI43/XI6/NET_001 XI31/XI1/XI43/NET36
+ XI31/XI1/XI43/XI6/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI6/MM_instance_269 XI31/XI1/XI43/XI6/NET_008
+ XI31/XI1/XI43/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_263 VDD! OP1<8> XI31/XI1/XI43/XI6/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI6/MM_instance_309 XI31/XI1/XI43/XI6/NET_011 OP1<8> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI6/MM_instance_297 VDD! XI31/XI1/XI43/NET36
+ XI31/XI1/XI43/XI6/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_303 XI31/XI1/XI43/XI6/NET_011
+ XI31/XI1/XI43/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_290 XI31/XI1/XI43/XI6/NET_005
+ XI31/XI1/XI43/XI6/NET_001 XI31/XI1/XI43/XI6/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_284 XI31/XI1/XI43/XI6/NET_010 XI31/XI1/XI43/NET36
+ XI31/XI1/XI43/XI6/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI6/MM_instance_280 XI31/XI1/XI43/XI6/NET_009 OP1<8>
+ XI31/XI1/XI43/XI6/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_275 VDD! XI31/XI1/XI43/OP0_TEMP<1>
+ XI31/XI1/XI43/XI6/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI6/MM_instance_315 XI31/XI1/XI43/S_1<1>
+ XI31/XI1/XI43/XI6/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI1/MM_instance_159 XI31/XI1/XI43/NET21 XI31/XI1/XI43/XI1/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI1/MM_instance_166 VSS! OP1<8> XI31/XI1/XI43/XI1/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_170 XI31/XI1/XI43/XI1/NET_000
+ XI31/XI1/XI43/OP0_TEMP<1> XI31/XI1/XI43/XI1/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_176 XI31/XI1/XI43/XI1/NET_001 XI31/XI1/XI43/NET16
+ XI31/XI1/XI43/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI1/MM_instance_188 XI31/XI1/XI43/XI1/NET_002
+ XI31/XI1/XI43/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_182 VSS! OP1<8> XI31/XI1/XI43/XI1/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI1/MM_instance_227 XI31/XI1/XI43/XI1/NET_006 OP1<8> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI1/MM_instance_215 VSS! XI31/XI1/XI43/NET16
+ XI31/XI1/XI43/XI1/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_221 XI31/XI1/XI43/XI1/NET_006
+ XI31/XI1/XI43/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_209 XI31/XI1/XI43/XI1/NET_005
+ XI31/XI1/XI43/XI1/NET_001 XI31/XI1/XI43/XI1/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_203 XI31/XI1/XI43/XI1/NET_004 XI31/XI1/XI43/NET16
+ XI31/XI1/XI43/XI1/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI1/MM_instance_199 XI31/XI1/XI43/XI1/NET_003 OP1<8>
+ XI31/XI1/XI43/XI1/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_194 VSS! XI31/XI1/XI43/OP0_TEMP<1>
+ XI31/XI1/XI43/XI1/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI1/MM_instance_233 XI31/XI1/XI43/S_0<1>
+ XI31/XI1/XI43/XI1/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI1/MM_instance_239 XI31/XI1/XI43/NET21 XI31/XI1/XI43/XI1/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI1/MM_instance_246 VDD! OP1<8> XI31/XI1/XI43/XI1/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_251 XI31/XI1/XI43/XI1/NET_007
+ XI31/XI1/XI43/OP0_TEMP<1> XI31/XI1/XI43/XI1/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_257 XI31/XI1/XI43/XI1/NET_001 XI31/XI1/XI43/NET16
+ XI31/XI1/XI43/XI1/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI1/MM_instance_269 XI31/XI1/XI43/XI1/NET_008
+ XI31/XI1/XI43/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_263 VDD! OP1<8> XI31/XI1/XI43/XI1/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI1/MM_instance_309 XI31/XI1/XI43/XI1/NET_011 OP1<8> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI1/MM_instance_297 VDD! XI31/XI1/XI43/NET16
+ XI31/XI1/XI43/XI1/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_303 XI31/XI1/XI43/XI1/NET_011
+ XI31/XI1/XI43/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_290 XI31/XI1/XI43/XI1/NET_005
+ XI31/XI1/XI43/XI1/NET_001 XI31/XI1/XI43/XI1/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_284 XI31/XI1/XI43/XI1/NET_010 XI31/XI1/XI43/NET16
+ XI31/XI1/XI43/XI1/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI1/MM_instance_280 XI31/XI1/XI43/XI1/NET_009 OP1<8>
+ XI31/XI1/XI43/XI1/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_275 VDD! XI31/XI1/XI43/OP0_TEMP<1>
+ XI31/XI1/XI43/XI1/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI1/MM_instance_315 XI31/XI1/XI43/S_0<1>
+ XI31/XI1/XI43/XI1/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI7/MM_instance_159 XI31/XI1/XI43/NET46 XI31/XI1/XI43/XI7/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI7/MM_instance_166 VSS! OP1<9> XI31/XI1/XI43/XI7/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_170 XI31/XI1/XI43/XI7/NET_000
+ XI31/XI1/XI43/OP0_TEMP<2> XI31/XI1/XI43/XI7/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_176 XI31/XI1/XI43/XI7/NET_001 XI31/XI1/XI43/NET41
+ XI31/XI1/XI43/XI7/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI7/MM_instance_188 XI31/XI1/XI43/XI7/NET_002
+ XI31/XI1/XI43/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_182 VSS! OP1<9> XI31/XI1/XI43/XI7/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI7/MM_instance_227 XI31/XI1/XI43/XI7/NET_006 OP1<9> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI7/MM_instance_215 VSS! XI31/XI1/XI43/NET41
+ XI31/XI1/XI43/XI7/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_221 XI31/XI1/XI43/XI7/NET_006
+ XI31/XI1/XI43/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_209 XI31/XI1/XI43/XI7/NET_005
+ XI31/XI1/XI43/XI7/NET_001 XI31/XI1/XI43/XI7/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_203 XI31/XI1/XI43/XI7/NET_004 XI31/XI1/XI43/NET41
+ XI31/XI1/XI43/XI7/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI7/MM_instance_199 XI31/XI1/XI43/XI7/NET_003 OP1<9>
+ XI31/XI1/XI43/XI7/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_194 VSS! XI31/XI1/XI43/OP0_TEMP<2>
+ XI31/XI1/XI43/XI7/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI7/MM_instance_233 XI31/XI1/XI43/S_1<2>
+ XI31/XI1/XI43/XI7/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI7/MM_instance_239 XI31/XI1/XI43/NET46 XI31/XI1/XI43/XI7/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI7/MM_instance_246 VDD! OP1<9> XI31/XI1/XI43/XI7/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_251 XI31/XI1/XI43/XI7/NET_007
+ XI31/XI1/XI43/OP0_TEMP<2> XI31/XI1/XI43/XI7/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_257 XI31/XI1/XI43/XI7/NET_001 XI31/XI1/XI43/NET41
+ XI31/XI1/XI43/XI7/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI7/MM_instance_269 XI31/XI1/XI43/XI7/NET_008
+ XI31/XI1/XI43/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_263 VDD! OP1<9> XI31/XI1/XI43/XI7/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI7/MM_instance_309 XI31/XI1/XI43/XI7/NET_011 OP1<9> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI7/MM_instance_297 VDD! XI31/XI1/XI43/NET41
+ XI31/XI1/XI43/XI7/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_303 XI31/XI1/XI43/XI7/NET_011
+ XI31/XI1/XI43/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_290 XI31/XI1/XI43/XI7/NET_005
+ XI31/XI1/XI43/XI7/NET_001 XI31/XI1/XI43/XI7/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_284 XI31/XI1/XI43/XI7/NET_010 XI31/XI1/XI43/NET41
+ XI31/XI1/XI43/XI7/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI7/MM_instance_280 XI31/XI1/XI43/XI7/NET_009 OP1<9>
+ XI31/XI1/XI43/XI7/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_275 VDD! XI31/XI1/XI43/OP0_TEMP<2>
+ XI31/XI1/XI43/XI7/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI7/MM_instance_315 XI31/XI1/XI43/S_1<2>
+ XI31/XI1/XI43/XI7/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI2/MM_instance_159 XI31/XI1/XI43/NET26 XI31/XI1/XI43/XI2/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI2/MM_instance_166 VSS! OP1<9> XI31/XI1/XI43/XI2/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_170 XI31/XI1/XI43/XI2/NET_000
+ XI31/XI1/XI43/OP0_TEMP<2> XI31/XI1/XI43/XI2/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_176 XI31/XI1/XI43/XI2/NET_001 XI31/XI1/XI43/NET21
+ XI31/XI1/XI43/XI2/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI2/MM_instance_188 XI31/XI1/XI43/XI2/NET_002
+ XI31/XI1/XI43/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_182 VSS! OP1<9> XI31/XI1/XI43/XI2/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI2/MM_instance_227 XI31/XI1/XI43/XI2/NET_006 OP1<9> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI2/MM_instance_215 VSS! XI31/XI1/XI43/NET21
+ XI31/XI1/XI43/XI2/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_221 XI31/XI1/XI43/XI2/NET_006
+ XI31/XI1/XI43/OP0_TEMP<2> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_209 XI31/XI1/XI43/XI2/NET_005
+ XI31/XI1/XI43/XI2/NET_001 XI31/XI1/XI43/XI2/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_203 XI31/XI1/XI43/XI2/NET_004 XI31/XI1/XI43/NET21
+ XI31/XI1/XI43/XI2/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI2/MM_instance_199 XI31/XI1/XI43/XI2/NET_003 OP1<9>
+ XI31/XI1/XI43/XI2/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_194 VSS! XI31/XI1/XI43/OP0_TEMP<2>
+ XI31/XI1/XI43/XI2/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI2/MM_instance_233 XI31/XI1/XI43/S_0<2>
+ XI31/XI1/XI43/XI2/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI2/MM_instance_239 XI31/XI1/XI43/NET26 XI31/XI1/XI43/XI2/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI2/MM_instance_246 VDD! OP1<9> XI31/XI1/XI43/XI2/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_251 XI31/XI1/XI43/XI2/NET_007
+ XI31/XI1/XI43/OP0_TEMP<2> XI31/XI1/XI43/XI2/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_257 XI31/XI1/XI43/XI2/NET_001 XI31/XI1/XI43/NET21
+ XI31/XI1/XI43/XI2/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI2/MM_instance_269 XI31/XI1/XI43/XI2/NET_008
+ XI31/XI1/XI43/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_263 VDD! OP1<9> XI31/XI1/XI43/XI2/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI2/MM_instance_309 XI31/XI1/XI43/XI2/NET_011 OP1<9> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI2/MM_instance_297 VDD! XI31/XI1/XI43/NET21
+ XI31/XI1/XI43/XI2/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_303 XI31/XI1/XI43/XI2/NET_011
+ XI31/XI1/XI43/OP0_TEMP<2> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_290 XI31/XI1/XI43/XI2/NET_005
+ XI31/XI1/XI43/XI2/NET_001 XI31/XI1/XI43/XI2/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_284 XI31/XI1/XI43/XI2/NET_010 XI31/XI1/XI43/NET21
+ XI31/XI1/XI43/XI2/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI2/MM_instance_280 XI31/XI1/XI43/XI2/NET_009 OP1<9>
+ XI31/XI1/XI43/XI2/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_275 VDD! XI31/XI1/XI43/OP0_TEMP<2>
+ XI31/XI1/XI43/XI2/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI2/MM_instance_315 XI31/XI1/XI43/S_0<2>
+ XI31/XI1/XI43/XI2/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI8/MM_instance_159 XI31/XI1/XI43/CO_1 XI31/XI1/XI43/XI8/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI8/MM_instance_166 VSS! OP1<10> XI31/XI1/XI43/XI8/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_170 XI31/XI1/XI43/XI8/NET_000 XI31/XI1/NET18
+ XI31/XI1/XI43/XI8/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_176 XI31/XI1/XI43/XI8/NET_001 XI31/XI1/XI43/NET46
+ XI31/XI1/XI43/XI8/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI8/MM_instance_188 XI31/XI1/XI43/XI8/NET_002 XI31/XI1/NET18 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_182 VSS! OP1<10> XI31/XI1/XI43/XI8/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI8/MM_instance_227 XI31/XI1/XI43/XI8/NET_006 OP1<10> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI8/MM_instance_215 VSS! XI31/XI1/XI43/NET46
+ XI31/XI1/XI43/XI8/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_221 XI31/XI1/XI43/XI8/NET_006 XI31/XI1/NET18 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_209 XI31/XI1/XI43/XI8/NET_005
+ XI31/XI1/XI43/XI8/NET_001 XI31/XI1/XI43/XI8/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_203 XI31/XI1/XI43/XI8/NET_004 XI31/XI1/XI43/NET46
+ XI31/XI1/XI43/XI8/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI8/MM_instance_199 XI31/XI1/XI43/XI8/NET_003 OP1<10>
+ XI31/XI1/XI43/XI8/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_194 VSS! XI31/XI1/NET18 XI31/XI1/XI43/XI8/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI8/MM_instance_233 XI31/XI1/XI43/S_1<3>
+ XI31/XI1/XI43/XI8/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI8/MM_instance_239 XI31/XI1/XI43/CO_1 XI31/XI1/XI43/XI8/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI8/MM_instance_246 VDD! OP1<10> XI31/XI1/XI43/XI8/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_251 XI31/XI1/XI43/XI8/NET_007 XI31/XI1/NET18
+ XI31/XI1/XI43/XI8/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_257 XI31/XI1/XI43/XI8/NET_001 XI31/XI1/XI43/NET46
+ XI31/XI1/XI43/XI8/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI8/MM_instance_269 XI31/XI1/XI43/XI8/NET_008 XI31/XI1/NET18 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_263 VDD! OP1<10> XI31/XI1/XI43/XI8/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI8/MM_instance_309 XI31/XI1/XI43/XI8/NET_011 OP1<10> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI8/MM_instance_297 VDD! XI31/XI1/XI43/NET46
+ XI31/XI1/XI43/XI8/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_303 XI31/XI1/XI43/XI8/NET_011 XI31/XI1/NET18 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_290 XI31/XI1/XI43/XI8/NET_005
+ XI31/XI1/XI43/XI8/NET_001 XI31/XI1/XI43/XI8/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_284 XI31/XI1/XI43/XI8/NET_010 XI31/XI1/XI43/NET46
+ XI31/XI1/XI43/XI8/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI8/MM_instance_280 XI31/XI1/XI43/XI8/NET_009 OP1<10>
+ XI31/XI1/XI43/XI8/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_275 VDD! XI31/XI1/NET18 XI31/XI1/XI43/XI8/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI8/MM_instance_315 XI31/XI1/XI43/S_1<3>
+ XI31/XI1/XI43/XI8/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI43/XI3/MM_instance_159 XI31/XI1/XI43/CO_0 XI31/XI1/XI43/XI3/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI43/XI3/MM_instance_166 VSS! OP1<10> XI31/XI1/XI43/XI3/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_170 XI31/XI1/XI43/XI3/NET_000 XI31/XI1/NET18
+ XI31/XI1/XI43/XI3/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_176 XI31/XI1/XI43/XI3/NET_001 XI31/XI1/XI43/NET26
+ XI31/XI1/XI43/XI3/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI43/XI3/MM_instance_188 XI31/XI1/XI43/XI3/NET_002 XI31/XI1/NET18 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_182 VSS! OP1<10> XI31/XI1/XI43/XI3/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI3/MM_instance_227 XI31/XI1/XI43/XI3/NET_006 OP1<10> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI43/XI3/MM_instance_215 VSS! XI31/XI1/XI43/NET26
+ XI31/XI1/XI43/XI3/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_221 XI31/XI1/XI43/XI3/NET_006 XI31/XI1/NET18 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_209 XI31/XI1/XI43/XI3/NET_005
+ XI31/XI1/XI43/XI3/NET_001 XI31/XI1/XI43/XI3/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_203 XI31/XI1/XI43/XI3/NET_004 XI31/XI1/XI43/NET26
+ XI31/XI1/XI43/XI3/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI43/XI3/MM_instance_199 XI31/XI1/XI43/XI3/NET_003 OP1<10>
+ XI31/XI1/XI43/XI3/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_194 VSS! XI31/XI1/NET18 XI31/XI1/XI43/XI3/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI43/XI3/MM_instance_233 XI31/XI1/XI43/S_0<3>
+ XI31/XI1/XI43/XI3/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI43/XI3/MM_instance_239 XI31/XI1/XI43/CO_0 XI31/XI1/XI43/XI3/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI43/XI3/MM_instance_246 VDD! OP1<10> XI31/XI1/XI43/XI3/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_251 XI31/XI1/XI43/XI3/NET_007 XI31/XI1/NET18
+ XI31/XI1/XI43/XI3/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_257 XI31/XI1/XI43/XI3/NET_001 XI31/XI1/XI43/NET26
+ XI31/XI1/XI43/XI3/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI43/XI3/MM_instance_269 XI31/XI1/XI43/XI3/NET_008 XI31/XI1/NET18 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_263 VDD! OP1<10> XI31/XI1/XI43/XI3/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI3/MM_instance_309 XI31/XI1/XI43/XI3/NET_011 OP1<10> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI43/XI3/MM_instance_297 VDD! XI31/XI1/XI43/NET26
+ XI31/XI1/XI43/XI3/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_303 XI31/XI1/XI43/XI3/NET_011 XI31/XI1/NET18 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_290 XI31/XI1/XI43/XI3/NET_005
+ XI31/XI1/XI43/XI3/NET_001 XI31/XI1/XI43/XI3/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_284 XI31/XI1/XI43/XI3/NET_010 XI31/XI1/XI43/NET26
+ XI31/XI1/XI43/XI3/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI43/XI3/MM_instance_280 XI31/XI1/XI43/XI3/NET_009 OP1<10>
+ XI31/XI1/XI43/XI3/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_275 VDD! XI31/XI1/NET18 XI31/XI1/XI43/XI3/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI43/XI3/MM_instance_315 XI31/XI1/XI43/S_0<3>
+ XI31/XI1/XI43/XI3/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI17/MM_i_10 VSS! XI31/XI1/NET3 XI31/XI1/XI42/XI17/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI17/MM_i_4 XI31/XI1/XI42/XI17/NET_1 XI31/XI1/XI42/S_0<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI17/MM_i_5 XI31/XI1/XI42/XI17/Z_NEG XI31/XI1/XI42/XI17/X1
+ XI31/XI1/XI42/XI17/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI17/MM_i_2 XI31/XI1/XI42/XI17/Z_NEG XI31/XI1/NET3
+ XI31/XI1/XI42/XI17/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI17/MM_i_3 XI31/XI1/XI42/XI17/NET_0 XI31/XI1/XI42/S_1<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI42/XI17/MM_i_0 XI31/ARITHMETIC_OUT<4> XI31/XI1/XI42/XI17/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI17/MM_i_11 VDD! XI31/XI1/NET3 XI31/XI1/XI42/XI17/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI17/MM_i_8 VDD! XI31/XI1/XI42/S_0<0> XI31/XI1/XI42/XI17/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI17/MM_i_6 XI31/XI1/XI42/XI17/NET_2 XI31/XI1/NET3
+ XI31/XI1/XI42/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI17/MM_i_9 XI31/XI1/XI42/XI17/NET_3 XI31/XI1/XI42/XI17/X1
+ XI31/XI1/XI42/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI17/MM_i_7 VDD! XI31/XI1/XI42/S_1<0> XI31/XI1/XI42/XI17/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI17/MM_i_1 XI31/ARITHMETIC_OUT<4> XI31/XI1/XI42/XI17/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI25/MM_i_10 VSS! XI31/XI1/NET3 XI31/XI1/XI42/XI25/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI25/MM_i_4 XI31/XI1/XI42/XI25/NET_1 XI31/XI1/XI42/S_0<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI25/MM_i_5 XI31/XI1/XI42/XI25/Z_NEG XI31/XI1/XI42/XI25/X1
+ XI31/XI1/XI42/XI25/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI25/MM_i_2 XI31/XI1/XI42/XI25/Z_NEG XI31/XI1/NET3
+ XI31/XI1/XI42/XI25/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI25/MM_i_3 XI31/XI1/XI42/XI25/NET_0 XI31/XI1/XI42/S_1<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI42/XI25/MM_i_0 XI31/ARITHMETIC_OUT<5> XI31/XI1/XI42/XI25/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI25/MM_i_11 VDD! XI31/XI1/NET3 XI31/XI1/XI42/XI25/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI25/MM_i_8 VDD! XI31/XI1/XI42/S_0<1> XI31/XI1/XI42/XI25/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI25/MM_i_6 XI31/XI1/XI42/XI25/NET_2 XI31/XI1/NET3
+ XI31/XI1/XI42/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI25/MM_i_9 XI31/XI1/XI42/XI25/NET_3 XI31/XI1/XI42/XI25/X1
+ XI31/XI1/XI42/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI25/MM_i_7 VDD! XI31/XI1/XI42/S_1<1> XI31/XI1/XI42/XI25/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI25/MM_i_1 XI31/ARITHMETIC_OUT<5> XI31/XI1/XI42/XI25/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI26/MM_i_10 VSS! XI31/XI1/NET3 XI31/XI1/XI42/XI26/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI26/MM_i_4 XI31/XI1/XI42/XI26/NET_1 XI31/XI1/XI42/S_0<2> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI26/MM_i_5 XI31/XI1/XI42/XI26/Z_NEG XI31/XI1/XI42/XI26/X1
+ XI31/XI1/XI42/XI26/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI26/MM_i_2 XI31/XI1/XI42/XI26/Z_NEG XI31/XI1/NET3
+ XI31/XI1/XI42/XI26/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI26/MM_i_3 XI31/XI1/XI42/XI26/NET_0 XI31/XI1/XI42/S_1<2> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI42/XI26/MM_i_0 XI31/ARITHMETIC_OUT<6> XI31/XI1/XI42/XI26/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI26/MM_i_11 VDD! XI31/XI1/NET3 XI31/XI1/XI42/XI26/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI26/MM_i_8 VDD! XI31/XI1/XI42/S_0<2> XI31/XI1/XI42/XI26/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI26/MM_i_6 XI31/XI1/XI42/XI26/NET_2 XI31/XI1/NET3
+ XI31/XI1/XI42/XI26/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI26/MM_i_9 XI31/XI1/XI42/XI26/NET_3 XI31/XI1/XI42/XI26/X1
+ XI31/XI1/XI42/XI26/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI26/MM_i_7 VDD! XI31/XI1/XI42/S_1<2> XI31/XI1/XI42/XI26/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI26/MM_i_1 XI31/ARITHMETIC_OUT<6> XI31/XI1/XI42/XI26/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI18/MM_i_10 VSS! XI31/XI1/NET3 XI31/XI1/XI42/XI18/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI18/MM_i_4 XI31/XI1/XI42/XI18/NET_1 XI31/XI1/XI42/CO_0 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI18/MM_i_5 XI31/XI1/XI42/XI18/Z_NEG XI31/XI1/XI42/XI18/X1
+ XI31/XI1/XI42/XI18/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI18/MM_i_2 XI31/XI1/XI42/XI18/Z_NEG XI31/XI1/NET3
+ XI31/XI1/XI42/XI18/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI18/MM_i_3 XI31/XI1/XI42/XI18/NET_0 XI31/XI1/XI42/CO_1 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI42/XI18/MM_i_0 XI31/XI1/NET12 XI31/XI1/XI42/XI18/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI18/MM_i_11 VDD! XI31/XI1/NET3 XI31/XI1/XI42/XI18/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI18/MM_i_8 VDD! XI31/XI1/XI42/CO_0 XI31/XI1/XI42/XI18/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI18/MM_i_6 XI31/XI1/XI42/XI18/NET_2 XI31/XI1/NET3
+ XI31/XI1/XI42/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI18/MM_i_9 XI31/XI1/XI42/XI18/NET_3 XI31/XI1/XI42/XI18/X1
+ XI31/XI1/XI42/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI18/MM_i_7 VDD! XI31/XI1/XI42/CO_1 XI31/XI1/XI42/XI18/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI18/MM_i_1 XI31/XI1/NET12 XI31/XI1/XI42/XI18/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI9/MM_i_0 XI31/XI1/XI42/XI9/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI9/MM_i_7 VSS! OP0<4> XI31/XI1/XI42/XI9/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI42/XI9/MM_i_13 XI31/XI1/XI42/OP0_TEMP<0> XI31/XI1/XI42/XI9/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI42/XI9/MM_i_19 XI31/XI1/XI42/XI9/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI42/OP0_TEMP<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI42/XI9/MM_i_24 VSS! OP0<4> XI31/XI1/XI42/XI9/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI9/MM_i_30 XI31/XI1/XI42/XI9/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI42/XI9/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI9/MM_i_35 VDD! OP0<4> XI31/XI1/XI42/XI9/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI42/XI9/MM_i_41 XI31/XI1/XI42/XI9/NET_003 XI31/XI1/XI42/XI9/NET_000
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI1/XI42/XI9/MM_i_47 XI31/XI1/XI42/OP0_TEMP<0> CTRL_BUFF<0>
+ XI31/XI1/XI42/XI9/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI42/XI9/MM_i_53 XI31/XI1/XI42/XI9/NET_003 OP0<4>
+ XI31/XI1/XI42/OP0_TEMP<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI10/MM_i_0 XI31/XI1/XI42/XI10/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI10/MM_i_7 VSS! OP0<5> XI31/XI1/XI42/XI10/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI42/XI10/MM_i_13 XI31/XI1/XI42/OP0_TEMP<1> XI31/XI1/XI42/XI10/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI42/XI10/MM_i_19 XI31/XI1/XI42/XI10/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI42/OP0_TEMP<1> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI42/XI10/MM_i_24 VSS! OP0<5> XI31/XI1/XI42/XI10/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI10/MM_i_30 XI31/XI1/XI42/XI10/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI42/XI10/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI10/MM_i_35 VDD! OP0<5> XI31/XI1/XI42/XI10/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI42/XI10/MM_i_41 XI31/XI1/XI42/XI10/NET_003
+ XI31/XI1/XI42/XI10/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI42/XI10/MM_i_47 XI31/XI1/XI42/OP0_TEMP<1> CTRL_BUFF<0>
+ XI31/XI1/XI42/XI10/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI42/XI10/MM_i_53 XI31/XI1/XI42/XI10/NET_003 OP0<5>
+ XI31/XI1/XI42/OP0_TEMP<1> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI11/MM_i_0 XI31/XI1/XI42/XI11/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI11/MM_i_7 VSS! OP0<6> XI31/XI1/XI42/XI11/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI42/XI11/MM_i_13 XI31/XI1/NET11 XI31/XI1/XI42/XI11/NET_000 VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06
mXI31/XI1/XI42/XI11/MM_i_19 XI31/XI1/XI42/XI11/NET_001 CTRL_BUFF<0>
+ XI31/XI1/NET11 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14
+ PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI42/XI11/MM_i_24 VSS! OP0<6> XI31/XI1/XI42/XI11/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI11/MM_i_30 XI31/XI1/XI42/XI11/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI42/XI11/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI11/MM_i_35 VDD! OP0<6> XI31/XI1/XI42/XI11/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI42/XI11/MM_i_41 XI31/XI1/XI42/XI11/NET_003
+ XI31/XI1/XI42/XI11/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI42/XI11/MM_i_47 XI31/XI1/NET11 CTRL_BUFF<0>
+ XI31/XI1/XI42/XI11/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI42/XI11/MM_i_53 XI31/XI1/XI42/XI11/NET_003 OP0<6> XI31/XI1/NET11
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI5/MM_instance_159 XI31/XI1/XI42/NET36 XI31/XI1/XI42/XI5/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI5/MM_instance_166 VSS! OP1<4> XI31/XI1/XI42/XI5/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_170 XI31/XI1/XI42/XI5/NET_000
+ XI31/XI1/XI42/OP0_TEMP<0> XI31/XI1/XI42/XI5/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_176 XI31/XI1/XI42/XI5/NET_001 VDD!
+ XI31/XI1/XI42/XI5/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI42/XI5/MM_instance_188 XI31/XI1/XI42/XI5/NET_002
+ XI31/XI1/XI42/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_182 VSS! OP1<4> XI31/XI1/XI42/XI5/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI5/MM_instance_227 XI31/XI1/XI42/XI5/NET_006 OP1<4> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI5/MM_instance_215 VSS! VDD! XI31/XI1/XI42/XI5/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_221 XI31/XI1/XI42/XI5/NET_006
+ XI31/XI1/XI42/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_209 XI31/XI1/XI42/XI5/NET_005
+ XI31/XI1/XI42/XI5/NET_001 XI31/XI1/XI42/XI5/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_203 XI31/XI1/XI42/XI5/NET_004 VDD!
+ XI31/XI1/XI42/XI5/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI42/XI5/MM_instance_199 XI31/XI1/XI42/XI5/NET_003 OP1<4>
+ XI31/XI1/XI42/XI5/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_194 VSS! XI31/XI1/XI42/OP0_TEMP<0>
+ XI31/XI1/XI42/XI5/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI5/MM_instance_233 XI31/XI1/XI42/S_1<0>
+ XI31/XI1/XI42/XI5/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI5/MM_instance_239 XI31/XI1/XI42/NET36 XI31/XI1/XI42/XI5/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI5/MM_instance_246 VDD! OP1<4> XI31/XI1/XI42/XI5/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_251 XI31/XI1/XI42/XI5/NET_007
+ XI31/XI1/XI42/OP0_TEMP<0> XI31/XI1/XI42/XI5/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_257 XI31/XI1/XI42/XI5/NET_001 VDD!
+ XI31/XI1/XI42/XI5/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI42/XI5/MM_instance_269 XI31/XI1/XI42/XI5/NET_008
+ XI31/XI1/XI42/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_263 VDD! OP1<4> XI31/XI1/XI42/XI5/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI5/MM_instance_309 XI31/XI1/XI42/XI5/NET_011 OP1<4> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI5/MM_instance_297 VDD! VDD! XI31/XI1/XI42/XI5/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_303 XI31/XI1/XI42/XI5/NET_011
+ XI31/XI1/XI42/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_290 XI31/XI1/XI42/XI5/NET_005
+ XI31/XI1/XI42/XI5/NET_001 XI31/XI1/XI42/XI5/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_284 XI31/XI1/XI42/XI5/NET_010 VDD!
+ XI31/XI1/XI42/XI5/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI42/XI5/MM_instance_280 XI31/XI1/XI42/XI5/NET_009 OP1<4>
+ XI31/XI1/XI42/XI5/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_275 VDD! XI31/XI1/XI42/OP0_TEMP<0>
+ XI31/XI1/XI42/XI5/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI5/MM_instance_315 XI31/XI1/XI42/S_1<0>
+ XI31/XI1/XI42/XI5/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI0/MM_instance_159 XI31/XI1/XI42/NET16 XI31/XI1/XI42/XI0/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI0/MM_instance_166 VSS! OP1<4> XI31/XI1/XI42/XI0/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_170 XI31/XI1/XI42/XI0/NET_000
+ XI31/XI1/XI42/OP0_TEMP<0> XI31/XI1/XI42/XI0/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_176 XI31/XI1/XI42/XI0/NET_001 VSS!
+ XI31/XI1/XI42/XI0/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI42/XI0/MM_instance_188 XI31/XI1/XI42/XI0/NET_002
+ XI31/XI1/XI42/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_182 VSS! OP1<4> XI31/XI1/XI42/XI0/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI0/MM_instance_227 XI31/XI1/XI42/XI0/NET_006 OP1<4> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI0/MM_instance_215 VSS! VSS! XI31/XI1/XI42/XI0/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_221 XI31/XI1/XI42/XI0/NET_006
+ XI31/XI1/XI42/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_209 XI31/XI1/XI42/XI0/NET_005
+ XI31/XI1/XI42/XI0/NET_001 XI31/XI1/XI42/XI0/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_203 XI31/XI1/XI42/XI0/NET_004 VSS!
+ XI31/XI1/XI42/XI0/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI42/XI0/MM_instance_199 XI31/XI1/XI42/XI0/NET_003 OP1<4>
+ XI31/XI1/XI42/XI0/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_194 VSS! XI31/XI1/XI42/OP0_TEMP<0>
+ XI31/XI1/XI42/XI0/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI0/MM_instance_233 XI31/XI1/XI42/S_0<0>
+ XI31/XI1/XI42/XI0/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI0/MM_instance_239 XI31/XI1/XI42/NET16 XI31/XI1/XI42/XI0/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI0/MM_instance_246 VDD! OP1<4> XI31/XI1/XI42/XI0/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_251 XI31/XI1/XI42/XI0/NET_007
+ XI31/XI1/XI42/OP0_TEMP<0> XI31/XI1/XI42/XI0/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_257 XI31/XI1/XI42/XI0/NET_001 VSS!
+ XI31/XI1/XI42/XI0/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI42/XI0/MM_instance_269 XI31/XI1/XI42/XI0/NET_008
+ XI31/XI1/XI42/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_263 VDD! OP1<4> XI31/XI1/XI42/XI0/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI0/MM_instance_309 XI31/XI1/XI42/XI0/NET_011 OP1<4> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI0/MM_instance_297 VDD! VSS! XI31/XI1/XI42/XI0/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_303 XI31/XI1/XI42/XI0/NET_011
+ XI31/XI1/XI42/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_290 XI31/XI1/XI42/XI0/NET_005
+ XI31/XI1/XI42/XI0/NET_001 XI31/XI1/XI42/XI0/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_284 XI31/XI1/XI42/XI0/NET_010 VSS!
+ XI31/XI1/XI42/XI0/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI42/XI0/MM_instance_280 XI31/XI1/XI42/XI0/NET_009 OP1<4>
+ XI31/XI1/XI42/XI0/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_275 VDD! XI31/XI1/XI42/OP0_TEMP<0>
+ XI31/XI1/XI42/XI0/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI0/MM_instance_315 XI31/XI1/XI42/S_0<0>
+ XI31/XI1/XI42/XI0/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI6/MM_instance_159 XI31/XI1/XI42/NET41 XI31/XI1/XI42/XI6/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI6/MM_instance_166 VSS! OP1<5> XI31/XI1/XI42/XI6/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_170 XI31/XI1/XI42/XI6/NET_000
+ XI31/XI1/XI42/OP0_TEMP<1> XI31/XI1/XI42/XI6/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_176 XI31/XI1/XI42/XI6/NET_001 XI31/XI1/XI42/NET36
+ XI31/XI1/XI42/XI6/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI42/XI6/MM_instance_188 XI31/XI1/XI42/XI6/NET_002
+ XI31/XI1/XI42/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_182 VSS! OP1<5> XI31/XI1/XI42/XI6/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI6/MM_instance_227 XI31/XI1/XI42/XI6/NET_006 OP1<5> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI6/MM_instance_215 VSS! XI31/XI1/XI42/NET36
+ XI31/XI1/XI42/XI6/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_221 XI31/XI1/XI42/XI6/NET_006
+ XI31/XI1/XI42/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_209 XI31/XI1/XI42/XI6/NET_005
+ XI31/XI1/XI42/XI6/NET_001 XI31/XI1/XI42/XI6/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_203 XI31/XI1/XI42/XI6/NET_004 XI31/XI1/XI42/NET36
+ XI31/XI1/XI42/XI6/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI42/XI6/MM_instance_199 XI31/XI1/XI42/XI6/NET_003 OP1<5>
+ XI31/XI1/XI42/XI6/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_194 VSS! XI31/XI1/XI42/OP0_TEMP<1>
+ XI31/XI1/XI42/XI6/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI6/MM_instance_233 XI31/XI1/XI42/S_1<1>
+ XI31/XI1/XI42/XI6/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI6/MM_instance_239 XI31/XI1/XI42/NET41 XI31/XI1/XI42/XI6/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI6/MM_instance_246 VDD! OP1<5> XI31/XI1/XI42/XI6/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_251 XI31/XI1/XI42/XI6/NET_007
+ XI31/XI1/XI42/OP0_TEMP<1> XI31/XI1/XI42/XI6/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_257 XI31/XI1/XI42/XI6/NET_001 XI31/XI1/XI42/NET36
+ XI31/XI1/XI42/XI6/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI42/XI6/MM_instance_269 XI31/XI1/XI42/XI6/NET_008
+ XI31/XI1/XI42/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_263 VDD! OP1<5> XI31/XI1/XI42/XI6/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI6/MM_instance_309 XI31/XI1/XI42/XI6/NET_011 OP1<5> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI6/MM_instance_297 VDD! XI31/XI1/XI42/NET36
+ XI31/XI1/XI42/XI6/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_303 XI31/XI1/XI42/XI6/NET_011
+ XI31/XI1/XI42/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_290 XI31/XI1/XI42/XI6/NET_005
+ XI31/XI1/XI42/XI6/NET_001 XI31/XI1/XI42/XI6/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_284 XI31/XI1/XI42/XI6/NET_010 XI31/XI1/XI42/NET36
+ XI31/XI1/XI42/XI6/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI42/XI6/MM_instance_280 XI31/XI1/XI42/XI6/NET_009 OP1<5>
+ XI31/XI1/XI42/XI6/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_275 VDD! XI31/XI1/XI42/OP0_TEMP<1>
+ XI31/XI1/XI42/XI6/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI6/MM_instance_315 XI31/XI1/XI42/S_1<1>
+ XI31/XI1/XI42/XI6/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI1/MM_instance_159 XI31/XI1/XI42/NET21 XI31/XI1/XI42/XI1/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI1/MM_instance_166 VSS! OP1<5> XI31/XI1/XI42/XI1/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_170 XI31/XI1/XI42/XI1/NET_000
+ XI31/XI1/XI42/OP0_TEMP<1> XI31/XI1/XI42/XI1/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_176 XI31/XI1/XI42/XI1/NET_001 XI31/XI1/XI42/NET16
+ XI31/XI1/XI42/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI42/XI1/MM_instance_188 XI31/XI1/XI42/XI1/NET_002
+ XI31/XI1/XI42/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_182 VSS! OP1<5> XI31/XI1/XI42/XI1/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI1/MM_instance_227 XI31/XI1/XI42/XI1/NET_006 OP1<5> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI1/MM_instance_215 VSS! XI31/XI1/XI42/NET16
+ XI31/XI1/XI42/XI1/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_221 XI31/XI1/XI42/XI1/NET_006
+ XI31/XI1/XI42/OP0_TEMP<1> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_209 XI31/XI1/XI42/XI1/NET_005
+ XI31/XI1/XI42/XI1/NET_001 XI31/XI1/XI42/XI1/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_203 XI31/XI1/XI42/XI1/NET_004 XI31/XI1/XI42/NET16
+ XI31/XI1/XI42/XI1/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI42/XI1/MM_instance_199 XI31/XI1/XI42/XI1/NET_003 OP1<5>
+ XI31/XI1/XI42/XI1/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_194 VSS! XI31/XI1/XI42/OP0_TEMP<1>
+ XI31/XI1/XI42/XI1/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI1/MM_instance_233 XI31/XI1/XI42/S_0<1>
+ XI31/XI1/XI42/XI1/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI1/MM_instance_239 XI31/XI1/XI42/NET21 XI31/XI1/XI42/XI1/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI1/MM_instance_246 VDD! OP1<5> XI31/XI1/XI42/XI1/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_251 XI31/XI1/XI42/XI1/NET_007
+ XI31/XI1/XI42/OP0_TEMP<1> XI31/XI1/XI42/XI1/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_257 XI31/XI1/XI42/XI1/NET_001 XI31/XI1/XI42/NET16
+ XI31/XI1/XI42/XI1/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI42/XI1/MM_instance_269 XI31/XI1/XI42/XI1/NET_008
+ XI31/XI1/XI42/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_263 VDD! OP1<5> XI31/XI1/XI42/XI1/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI1/MM_instance_309 XI31/XI1/XI42/XI1/NET_011 OP1<5> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI1/MM_instance_297 VDD! XI31/XI1/XI42/NET16
+ XI31/XI1/XI42/XI1/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_303 XI31/XI1/XI42/XI1/NET_011
+ XI31/XI1/XI42/OP0_TEMP<1> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_290 XI31/XI1/XI42/XI1/NET_005
+ XI31/XI1/XI42/XI1/NET_001 XI31/XI1/XI42/XI1/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_284 XI31/XI1/XI42/XI1/NET_010 XI31/XI1/XI42/NET16
+ XI31/XI1/XI42/XI1/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI42/XI1/MM_instance_280 XI31/XI1/XI42/XI1/NET_009 OP1<5>
+ XI31/XI1/XI42/XI1/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_275 VDD! XI31/XI1/XI42/OP0_TEMP<1>
+ XI31/XI1/XI42/XI1/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI1/MM_instance_315 XI31/XI1/XI42/S_0<1>
+ XI31/XI1/XI42/XI1/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI7/MM_instance_159 XI31/XI1/XI42/CO_1 XI31/XI1/XI42/XI7/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI7/MM_instance_166 VSS! OP1<6> XI31/XI1/XI42/XI7/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_170 XI31/XI1/XI42/XI7/NET_000 XI31/XI1/NET11
+ XI31/XI1/XI42/XI7/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_176 XI31/XI1/XI42/XI7/NET_001 XI31/XI1/XI42/NET41
+ XI31/XI1/XI42/XI7/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI42/XI7/MM_instance_188 XI31/XI1/XI42/XI7/NET_002 XI31/XI1/NET11 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_182 VSS! OP1<6> XI31/XI1/XI42/XI7/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI7/MM_instance_227 XI31/XI1/XI42/XI7/NET_006 OP1<6> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI7/MM_instance_215 VSS! XI31/XI1/XI42/NET41
+ XI31/XI1/XI42/XI7/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_221 XI31/XI1/XI42/XI7/NET_006 XI31/XI1/NET11 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_209 XI31/XI1/XI42/XI7/NET_005
+ XI31/XI1/XI42/XI7/NET_001 XI31/XI1/XI42/XI7/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_203 XI31/XI1/XI42/XI7/NET_004 XI31/XI1/XI42/NET41
+ XI31/XI1/XI42/XI7/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI42/XI7/MM_instance_199 XI31/XI1/XI42/XI7/NET_003 OP1<6>
+ XI31/XI1/XI42/XI7/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_194 VSS! XI31/XI1/NET11 XI31/XI1/XI42/XI7/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI7/MM_instance_233 XI31/XI1/XI42/S_1<2>
+ XI31/XI1/XI42/XI7/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI7/MM_instance_239 XI31/XI1/XI42/CO_1 XI31/XI1/XI42/XI7/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI7/MM_instance_246 VDD! OP1<6> XI31/XI1/XI42/XI7/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_251 XI31/XI1/XI42/XI7/NET_007 XI31/XI1/NET11
+ XI31/XI1/XI42/XI7/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_257 XI31/XI1/XI42/XI7/NET_001 XI31/XI1/XI42/NET41
+ XI31/XI1/XI42/XI7/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI42/XI7/MM_instance_269 XI31/XI1/XI42/XI7/NET_008 XI31/XI1/NET11 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_263 VDD! OP1<6> XI31/XI1/XI42/XI7/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI7/MM_instance_309 XI31/XI1/XI42/XI7/NET_011 OP1<6> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI7/MM_instance_297 VDD! XI31/XI1/XI42/NET41
+ XI31/XI1/XI42/XI7/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_303 XI31/XI1/XI42/XI7/NET_011 XI31/XI1/NET11 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_290 XI31/XI1/XI42/XI7/NET_005
+ XI31/XI1/XI42/XI7/NET_001 XI31/XI1/XI42/XI7/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_284 XI31/XI1/XI42/XI7/NET_010 XI31/XI1/XI42/NET41
+ XI31/XI1/XI42/XI7/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI42/XI7/MM_instance_280 XI31/XI1/XI42/XI7/NET_009 OP1<6>
+ XI31/XI1/XI42/XI7/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_275 VDD! XI31/XI1/NET11 XI31/XI1/XI42/XI7/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI7/MM_instance_315 XI31/XI1/XI42/S_1<2>
+ XI31/XI1/XI42/XI7/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI42/XI2/MM_instance_159 XI31/XI1/XI42/CO_0 XI31/XI1/XI42/XI2/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI42/XI2/MM_instance_166 VSS! OP1<6> XI31/XI1/XI42/XI2/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_170 XI31/XI1/XI42/XI2/NET_000 XI31/XI1/NET11
+ XI31/XI1/XI42/XI2/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_176 XI31/XI1/XI42/XI2/NET_001 XI31/XI1/XI42/NET21
+ XI31/XI1/XI42/XI2/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI42/XI2/MM_instance_188 XI31/XI1/XI42/XI2/NET_002 XI31/XI1/NET11 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_182 VSS! OP1<6> XI31/XI1/XI42/XI2/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI2/MM_instance_227 XI31/XI1/XI42/XI2/NET_006 OP1<6> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI42/XI2/MM_instance_215 VSS! XI31/XI1/XI42/NET21
+ XI31/XI1/XI42/XI2/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_221 XI31/XI1/XI42/XI2/NET_006 XI31/XI1/NET11 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_209 XI31/XI1/XI42/XI2/NET_005
+ XI31/XI1/XI42/XI2/NET_001 XI31/XI1/XI42/XI2/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_203 XI31/XI1/XI42/XI2/NET_004 XI31/XI1/XI42/NET21
+ XI31/XI1/XI42/XI2/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI42/XI2/MM_instance_199 XI31/XI1/XI42/XI2/NET_003 OP1<6>
+ XI31/XI1/XI42/XI2/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_194 VSS! XI31/XI1/NET11 XI31/XI1/XI42/XI2/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI42/XI2/MM_instance_233 XI31/XI1/XI42/S_0<2>
+ XI31/XI1/XI42/XI2/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI42/XI2/MM_instance_239 XI31/XI1/XI42/CO_0 XI31/XI1/XI42/XI2/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI42/XI2/MM_instance_246 VDD! OP1<6> XI31/XI1/XI42/XI2/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_251 XI31/XI1/XI42/XI2/NET_007 XI31/XI1/NET11
+ XI31/XI1/XI42/XI2/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_257 XI31/XI1/XI42/XI2/NET_001 XI31/XI1/XI42/NET21
+ XI31/XI1/XI42/XI2/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI42/XI2/MM_instance_269 XI31/XI1/XI42/XI2/NET_008 XI31/XI1/NET11 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_263 VDD! OP1<6> XI31/XI1/XI42/XI2/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI2/MM_instance_309 XI31/XI1/XI42/XI2/NET_011 OP1<6> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI42/XI2/MM_instance_297 VDD! XI31/XI1/XI42/NET21
+ XI31/XI1/XI42/XI2/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_303 XI31/XI1/XI42/XI2/NET_011 XI31/XI1/NET11 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_290 XI31/XI1/XI42/XI2/NET_005
+ XI31/XI1/XI42/XI2/NET_001 XI31/XI1/XI42/XI2/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_284 XI31/XI1/XI42/XI2/NET_010 XI31/XI1/XI42/NET21
+ XI31/XI1/XI42/XI2/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI42/XI2/MM_instance_280 XI31/XI1/XI42/XI2/NET_009 OP1<6>
+ XI31/XI1/XI42/XI2/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_275 VDD! XI31/XI1/NET11 XI31/XI1/XI42/XI2/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI42/XI2/MM_instance_315 XI31/XI1/XI42/S_0<2>
+ XI31/XI1/XI42/XI2/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI17/MM_i_10 VSS! XI31/XI1/NET1 XI31/XI1/XI41/XI17/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI17/MM_i_4 XI31/XI1/XI41/XI17/NET_1 XI31/XI1/XI41/S_0<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI17/MM_i_5 XI31/XI1/XI41/XI17/Z_NEG XI31/XI1/XI41/XI17/X1
+ XI31/XI1/XI41/XI17/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI17/MM_i_2 XI31/XI1/XI41/XI17/Z_NEG XI31/XI1/NET1
+ XI31/XI1/XI41/XI17/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI17/MM_i_3 XI31/XI1/XI41/XI17/NET_0 XI31/XI1/XI41/S_1<0> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI41/XI17/MM_i_0 XI31/ARITHMETIC_OUT<2> XI31/XI1/XI41/XI17/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI41/XI17/MM_i_11 VDD! XI31/XI1/NET1 XI31/XI1/XI41/XI17/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI17/MM_i_8 VDD! XI31/XI1/XI41/S_0<0> XI31/XI1/XI41/XI17/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI17/MM_i_6 XI31/XI1/XI41/XI17/NET_2 XI31/XI1/NET1
+ XI31/XI1/XI41/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI17/MM_i_9 XI31/XI1/XI41/XI17/NET_3 XI31/XI1/XI41/XI17/X1
+ XI31/XI1/XI41/XI17/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI17/MM_i_7 VDD! XI31/XI1/XI41/S_1<0> XI31/XI1/XI41/XI17/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI41/XI17/MM_i_1 XI31/ARITHMETIC_OUT<2> XI31/XI1/XI41/XI17/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI41/XI25/MM_i_10 VSS! XI31/XI1/NET1 XI31/XI1/XI41/XI25/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI25/MM_i_4 XI31/XI1/XI41/XI25/NET_1 XI31/XI1/XI41/S_0<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI25/MM_i_5 XI31/XI1/XI41/XI25/Z_NEG XI31/XI1/XI41/XI25/X1
+ XI31/XI1/XI41/XI25/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI25/MM_i_2 XI31/XI1/XI41/XI25/Z_NEG XI31/XI1/NET1
+ XI31/XI1/XI41/XI25/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI25/MM_i_3 XI31/XI1/XI41/XI25/NET_0 XI31/XI1/XI41/S_1<1> VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI41/XI25/MM_i_0 XI31/ARITHMETIC_OUT<3> XI31/XI1/XI41/XI25/Z_NEG VSS!
+ VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI41/XI25/MM_i_11 VDD! XI31/XI1/NET1 XI31/XI1/XI41/XI25/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI25/MM_i_8 VDD! XI31/XI1/XI41/S_0<1> XI31/XI1/XI41/XI25/NET_2
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI25/MM_i_6 XI31/XI1/XI41/XI25/NET_2 XI31/XI1/NET1
+ XI31/XI1/XI41/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI25/MM_i_9 XI31/XI1/XI41/XI25/NET_3 XI31/XI1/XI41/XI25/X1
+ XI31/XI1/XI41/XI25/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI25/MM_i_7 VDD! XI31/XI1/XI41/S_1<1> XI31/XI1/XI41/XI25/NET_3
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI41/XI25/MM_i_1 XI31/ARITHMETIC_OUT<3> XI31/XI1/XI41/XI25/Z_NEG VDD!
+ VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI41/XI18/MM_i_10 VSS! XI31/XI1/NET1 XI31/XI1/XI41/XI18/X1 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI18/MM_i_4 XI31/XI1/XI41/XI18/NET_1 XI31/XI1/XI41/CO_0 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI18/MM_i_5 XI31/XI1/XI41/XI18/Z_NEG XI31/XI1/XI41/XI18/X1
+ XI31/XI1/XI41/XI18/NET_1 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI18/MM_i_2 XI31/XI1/XI41/XI18/Z_NEG XI31/XI1/NET1
+ XI31/XI1/XI41/XI18/NET_0 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI18/MM_i_3 XI31/XI1/XI41/XI18/NET_0 XI31/XI1/XI41/CO_1 VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06
mXI31/XI1/XI41/XI18/MM_i_0 XI31/XI1/NET3 XI31/XI1/XI41/XI18/Z_NEG VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI18/MM_i_11 VDD! XI31/XI1/NET1 XI31/XI1/XI41/XI18/X1 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI18/MM_i_8 VDD! XI31/XI1/XI41/CO_0 XI31/XI1/XI41/XI18/NET_2 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI18/MM_i_6 XI31/XI1/XI41/XI18/NET_2 XI31/XI1/NET1
+ XI31/XI1/XI41/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI18/MM_i_9 XI31/XI1/XI41/XI18/NET_3 XI31/XI1/XI41/XI18/X1
+ XI31/XI1/XI41/XI18/Z_NEG VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI18/MM_i_7 VDD! XI31/XI1/XI41/CO_1 XI31/XI1/XI41/XI18/NET_3 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI18/MM_i_1 XI31/XI1/NET3 XI31/XI1/XI41/XI18/Z_NEG VDD! VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI9/MM_i_0 XI31/XI1/XI41/XI9/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI9/MM_i_7 VSS! OP0<2> XI31/XI1/XI41/XI9/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI41/XI9/MM_i_13 XI31/XI1/XI41/OP0_TEMP<0> XI31/XI1/XI41/XI9/NET_000
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06
+ PS=1.12e-06
mXI31/XI1/XI41/XI9/MM_i_19 XI31/XI1/XI41/XI9/NET_001 CTRL_BUFF<0>
+ XI31/XI1/XI41/OP0_TEMP<0> VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14
+ AS=5.81e-14 PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI41/XI9/MM_i_24 VSS! OP0<2> XI31/XI1/XI41/XI9/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI9/MM_i_30 XI31/XI1/XI41/XI9/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI41/XI9/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI9/MM_i_35 VDD! OP0<2> XI31/XI1/XI41/XI9/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI41/XI9/MM_i_41 XI31/XI1/XI41/XI9/NET_003 XI31/XI1/XI41/XI9/NET_000
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06
+ PS=1.55e-06
mXI31/XI1/XI41/XI9/MM_i_47 XI31/XI1/XI41/OP0_TEMP<0> CTRL_BUFF<0>
+ XI31/XI1/XI41/XI9/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI41/XI9/MM_i_53 XI31/XI1/XI41/XI9/NET_003 OP0<2>
+ XI31/XI1/XI41/OP0_TEMP<0> VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI10/MM_i_0 XI31/XI1/XI41/XI10/NET_000 CTRL_BUFF<0> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI10/MM_i_7 VSS! OP0<3> XI31/XI1/XI41/XI10/NET_000 VSS! NMOS_VTL
+ L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07
mXI31/XI1/XI41/XI10/MM_i_13 XI31/XI1/NET2 XI31/XI1/XI41/XI10/NET_000 VSS! VSS!
+ NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06
mXI31/XI1/XI41/XI10/MM_i_19 XI31/XI1/XI41/XI10/NET_001 CTRL_BUFF<0>
+ XI31/XI1/NET2 VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14
+ PD=1.11e-06 PS=1.11e-06
mXI31/XI1/XI41/XI10/MM_i_24 VSS! OP0<3> XI31/XI1/XI41/XI10/NET_001 VSS! NMOS_VTL
+ L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI10/MM_i_30 XI31/XI1/XI41/XI10/NET_002 CTRL_BUFF<0>
+ XI31/XI1/XI41/XI10/NET_000 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI10/MM_i_35 VDD! OP0<3> XI31/XI1/XI41/XI10/NET_002 VDD! PMOS_VTL
+ L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07
mXI31/XI1/XI41/XI10/MM_i_41 XI31/XI1/XI41/XI10/NET_003
+ XI31/XI1/XI41/XI10/NET_000 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06
mXI31/XI1/XI41/XI10/MM_i_47 XI31/XI1/NET2 CTRL_BUFF<0>
+ XI31/XI1/XI41/XI10/NET_003 VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14
+ AS=8.82e-14 PD=1.54e-06 PS=1.54e-06
mXI31/XI1/XI41/XI10/MM_i_53 XI31/XI1/XI41/XI10/NET_003 OP0<3> XI31/XI1/NET2 VDD!
+ PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI5/MM_instance_159 XI31/XI1/XI41/NET36 XI31/XI1/XI41/XI5/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI41/XI5/MM_instance_166 VSS! OP1<2> XI31/XI1/XI41/XI5/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_170 XI31/XI1/XI41/XI5/NET_000
+ XI31/XI1/XI41/OP0_TEMP<0> XI31/XI1/XI41/XI5/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_176 XI31/XI1/XI41/XI5/NET_001 VDD!
+ XI31/XI1/XI41/XI5/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI41/XI5/MM_instance_188 XI31/XI1/XI41/XI5/NET_002
+ XI31/XI1/XI41/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_182 VSS! OP1<2> XI31/XI1/XI41/XI5/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI5/MM_instance_227 XI31/XI1/XI41/XI5/NET_006 OP1<2> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI5/MM_instance_215 VSS! VDD! XI31/XI1/XI41/XI5/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_221 XI31/XI1/XI41/XI5/NET_006
+ XI31/XI1/XI41/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_209 XI31/XI1/XI41/XI5/NET_005
+ XI31/XI1/XI41/XI5/NET_001 XI31/XI1/XI41/XI5/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_203 XI31/XI1/XI41/XI5/NET_004 VDD!
+ XI31/XI1/XI41/XI5/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI41/XI5/MM_instance_199 XI31/XI1/XI41/XI5/NET_003 OP1<2>
+ XI31/XI1/XI41/XI5/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_194 VSS! XI31/XI1/XI41/OP0_TEMP<0>
+ XI31/XI1/XI41/XI5/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI5/MM_instance_233 XI31/XI1/XI41/S_1<0>
+ XI31/XI1/XI41/XI5/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI5/MM_instance_239 XI31/XI1/XI41/NET36 XI31/XI1/XI41/XI5/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI41/XI5/MM_instance_246 VDD! OP1<2> XI31/XI1/XI41/XI5/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_251 XI31/XI1/XI41/XI5/NET_007
+ XI31/XI1/XI41/OP0_TEMP<0> XI31/XI1/XI41/XI5/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_257 XI31/XI1/XI41/XI5/NET_001 VDD!
+ XI31/XI1/XI41/XI5/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI41/XI5/MM_instance_269 XI31/XI1/XI41/XI5/NET_008
+ XI31/XI1/XI41/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_263 VDD! OP1<2> XI31/XI1/XI41/XI5/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI5/MM_instance_309 XI31/XI1/XI41/XI5/NET_011 OP1<2> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI5/MM_instance_297 VDD! VDD! XI31/XI1/XI41/XI5/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_303 XI31/XI1/XI41/XI5/NET_011
+ XI31/XI1/XI41/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_290 XI31/XI1/XI41/XI5/NET_005
+ XI31/XI1/XI41/XI5/NET_001 XI31/XI1/XI41/XI5/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_284 XI31/XI1/XI41/XI5/NET_010 VDD!
+ XI31/XI1/XI41/XI5/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI41/XI5/MM_instance_280 XI31/XI1/XI41/XI5/NET_009 OP1<2>
+ XI31/XI1/XI41/XI5/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_275 VDD! XI31/XI1/XI41/OP0_TEMP<0>
+ XI31/XI1/XI41/XI5/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI5/MM_instance_315 XI31/XI1/XI41/S_1<0>
+ XI31/XI1/XI41/XI5/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI0/MM_instance_159 XI31/XI1/XI41/NET16 XI31/XI1/XI41/XI0/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI41/XI0/MM_instance_166 VSS! OP1<2> XI31/XI1/XI41/XI0/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_170 XI31/XI1/XI41/XI0/NET_000
+ XI31/XI1/XI41/OP0_TEMP<0> XI31/XI1/XI41/XI0/NET_001 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_176 XI31/XI1/XI41/XI0/NET_001 VSS!
+ XI31/XI1/XI41/XI0/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI41/XI0/MM_instance_188 XI31/XI1/XI41/XI0/NET_002
+ XI31/XI1/XI41/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14
+ AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_182 VSS! OP1<2> XI31/XI1/XI41/XI0/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI0/MM_instance_227 XI31/XI1/XI41/XI0/NET_006 OP1<2> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI0/MM_instance_215 VSS! VSS! XI31/XI1/XI41/XI0/NET_006 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_221 XI31/XI1/XI41/XI0/NET_006
+ XI31/XI1/XI41/OP0_TEMP<0> VSS! VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_209 XI31/XI1/XI41/XI0/NET_005
+ XI31/XI1/XI41/XI0/NET_001 XI31/XI1/XI41/XI0/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_203 XI31/XI1/XI41/XI0/NET_004 VSS!
+ XI31/XI1/XI41/XI0/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI41/XI0/MM_instance_199 XI31/XI1/XI41/XI0/NET_003 OP1<2>
+ XI31/XI1/XI41/XI0/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_194 VSS! XI31/XI1/XI41/OP0_TEMP<0>
+ XI31/XI1/XI41/XI0/NET_003 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14
+ AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI0/MM_instance_233 XI31/XI1/XI41/S_0<0>
+ XI31/XI1/XI41/XI0/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI0/MM_instance_239 XI31/XI1/XI41/NET16 XI31/XI1/XI41/XI0/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI41/XI0/MM_instance_246 VDD! OP1<2> XI31/XI1/XI41/XI0/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_251 XI31/XI1/XI41/XI0/NET_007
+ XI31/XI1/XI41/OP0_TEMP<0> XI31/XI1/XI41/XI0/NET_001 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_257 XI31/XI1/XI41/XI0/NET_001 VSS!
+ XI31/XI1/XI41/XI0/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI41/XI0/MM_instance_269 XI31/XI1/XI41/XI0/NET_008
+ XI31/XI1/XI41/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14
+ AS=4.41e-14 PD=1.07e-06 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_263 VDD! OP1<2> XI31/XI1/XI41/XI0/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI0/MM_instance_309 XI31/XI1/XI41/XI0/NET_011 OP1<2> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI0/MM_instance_297 VDD! VSS! XI31/XI1/XI41/XI0/NET_011 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_303 XI31/XI1/XI41/XI0/NET_011
+ XI31/XI1/XI41/OP0_TEMP<0> VDD! VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_290 XI31/XI1/XI41/XI0/NET_005
+ XI31/XI1/XI41/XI0/NET_001 XI31/XI1/XI41/XI0/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_284 XI31/XI1/XI41/XI0/NET_010 VSS!
+ XI31/XI1/XI41/XI0/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI41/XI0/MM_instance_280 XI31/XI1/XI41/XI0/NET_009 OP1<2>
+ XI31/XI1/XI41/XI0/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_275 VDD! XI31/XI1/XI41/OP0_TEMP<0>
+ XI31/XI1/XI41/XI0/NET_009 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14
+ AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI0/MM_instance_315 XI31/XI1/XI41/S_0<0>
+ XI31/XI1/XI41/XI0/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI6/MM_instance_159 XI31/XI1/XI41/CO_1 XI31/XI1/XI41/XI6/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI41/XI6/MM_instance_166 VSS! OP1<3> XI31/XI1/XI41/XI6/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_170 XI31/XI1/XI41/XI6/NET_000 XI31/XI1/NET2
+ XI31/XI1/XI41/XI6/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_176 XI31/XI1/XI41/XI6/NET_001 XI31/XI1/XI41/NET36
+ XI31/XI1/XI41/XI6/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI41/XI6/MM_instance_188 XI31/XI1/XI41/XI6/NET_002 XI31/XI1/NET2 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_182 VSS! OP1<3> XI31/XI1/XI41/XI6/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI6/MM_instance_227 XI31/XI1/XI41/XI6/NET_006 OP1<3> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI6/MM_instance_215 VSS! XI31/XI1/XI41/NET36
+ XI31/XI1/XI41/XI6/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_221 XI31/XI1/XI41/XI6/NET_006 XI31/XI1/NET2 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_209 XI31/XI1/XI41/XI6/NET_005
+ XI31/XI1/XI41/XI6/NET_001 XI31/XI1/XI41/XI6/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_203 XI31/XI1/XI41/XI6/NET_004 XI31/XI1/XI41/NET36
+ XI31/XI1/XI41/XI6/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI41/XI6/MM_instance_199 XI31/XI1/XI41/XI6/NET_003 OP1<3>
+ XI31/XI1/XI41/XI6/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_194 VSS! XI31/XI1/NET2 XI31/XI1/XI41/XI6/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI6/MM_instance_233 XI31/XI1/XI41/S_1<1>
+ XI31/XI1/XI41/XI6/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI6/MM_instance_239 XI31/XI1/XI41/CO_1 XI31/XI1/XI41/XI6/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI41/XI6/MM_instance_246 VDD! OP1<3> XI31/XI1/XI41/XI6/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_251 XI31/XI1/XI41/XI6/NET_007 XI31/XI1/NET2
+ XI31/XI1/XI41/XI6/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_257 XI31/XI1/XI41/XI6/NET_001 XI31/XI1/XI41/NET36
+ XI31/XI1/XI41/XI6/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI41/XI6/MM_instance_269 XI31/XI1/XI41/XI6/NET_008 XI31/XI1/NET2 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_263 VDD! OP1<3> XI31/XI1/XI41/XI6/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI6/MM_instance_309 XI31/XI1/XI41/XI6/NET_011 OP1<3> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI6/MM_instance_297 VDD! XI31/XI1/XI41/NET36
+ XI31/XI1/XI41/XI6/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_303 XI31/XI1/XI41/XI6/NET_011 XI31/XI1/NET2 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_290 XI31/XI1/XI41/XI6/NET_005
+ XI31/XI1/XI41/XI6/NET_001 XI31/XI1/XI41/XI6/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_284 XI31/XI1/XI41/XI6/NET_010 XI31/XI1/XI41/NET36
+ XI31/XI1/XI41/XI6/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI41/XI6/MM_instance_280 XI31/XI1/XI41/XI6/NET_009 OP1<3>
+ XI31/XI1/XI41/XI6/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_275 VDD! XI31/XI1/NET2 XI31/XI1/XI41/XI6/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI41/XI6/MM_instance_315 XI31/XI1/XI41/S_1<1>
+ XI31/XI1/XI41/XI6/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
mXI31/XI1/XI41/XI1/MM_instance_159 XI31/XI1/XI41/CO_0 XI31/XI1/XI41/XI1/NET_001
+ VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06
+ PS=1.11e-06
mXI31/XI1/XI41/XI1/MM_instance_166 VSS! OP1<3> XI31/XI1/XI41/XI1/NET_000 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_170 XI31/XI1/XI41/XI1/NET_000 XI31/XI1/NET2
+ XI31/XI1/XI41/XI1/NET_001 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_176 XI31/XI1/XI41/XI1/NET_001 XI31/XI1/XI41/NET16
+ XI31/XI1/XI41/XI1/NET_002 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.045e-14 PD=7e-07 PS=7.1e-07
mXI31/XI1/XI41/XI1/MM_instance_188 XI31/XI1/XI41/XI1/NET_002 XI31/XI1/NET2 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_182 VSS! OP1<3> XI31/XI1/XI41/XI1/NET_002 VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI1/MM_instance_227 XI31/XI1/XI41/XI1/NET_006 OP1<3> VSS! VSS!
+ NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07
mXI31/XI1/XI41/XI1/MM_instance_215 VSS! XI31/XI1/XI41/NET16
+ XI31/XI1/XI41/XI1/NET_006 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_221 XI31/XI1/XI41/XI1/NET_006 XI31/XI1/NET2 VSS!
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_209 XI31/XI1/XI41/XI1/NET_005
+ XI31/XI1/XI41/XI1/NET_001 XI31/XI1/XI41/XI1/NET_006 VSS! NMOS_VTL L=5e-08
+ W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_203 XI31/XI1/XI41/XI1/NET_004 XI31/XI1/XI41/NET16
+ XI31/XI1/XI41/XI1/NET_005 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=3.15e-14 PD=7e-07 PS=7.2e-07
mXI31/XI1/XI41/XI1/MM_instance_199 XI31/XI1/XI41/XI1/NET_003 OP1<3>
+ XI31/XI1/XI41/XI1/NET_004 VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7e-07 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_194 VSS! XI31/XI1/NET2 XI31/XI1/XI41/XI1/NET_003
+ VSS! NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07
mXI31/XI1/XI41/XI1/MM_instance_233 XI31/XI1/XI41/S_0<1>
+ XI31/XI1/XI41/XI1/NET_005 VSS! VSS! NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14
+ AS=4.375e-14 PD=1.04e-06 PS=1.11e-06
mXI31/XI1/XI41/XI1/MM_instance_239 XI31/XI1/XI41/CO_0 XI31/XI1/XI41/XI1/NET_001
+ VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06
+ PS=1.54e-06
mXI31/XI1/XI41/XI1/MM_instance_246 VDD! OP1<3> XI31/XI1/XI41/XI1/NET_007 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_251 XI31/XI1/XI41/XI1/NET_007 XI31/XI1/NET2
+ XI31/XI1/XI41/XI1/NET_001 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_257 XI31/XI1/XI41/XI1/NET_001 XI31/XI1/XI41/NET16
+ XI31/XI1/XI41/XI1/NET_008 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.53e-14 PD=9.1e-07 PS=1.07e-06
mXI31/XI1/XI41/XI1/MM_instance_269 XI31/XI1/XI41/XI1/NET_008 XI31/XI1/NET2 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06
+ PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_263 VDD! OP1<3> XI31/XI1/XI41/XI1/NET_008 VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI1/MM_instance_309 XI31/XI1/XI41/XI1/NET_011 OP1<3> VDD! VDD!
+ PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07
mXI31/XI1/XI41/XI1/MM_instance_297 VDD! XI31/XI1/XI41/NET16
+ XI31/XI1/XI41/XI1/NET_011 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_303 XI31/XI1/XI41/XI1/NET_011 XI31/XI1/NET2 VDD!
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_290 XI31/XI1/XI41/XI1/NET_005
+ XI31/XI1/XI41/XI1/NET_001 XI31/XI1/XI41/XI1/NET_011 VDD! PMOS_VTL L=5e-08
+ W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_284 XI31/XI1/XI41/XI1/NET_010 XI31/XI1/XI41/NET16
+ XI31/XI1/XI41/XI1/NET_005 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.725e-14 PD=9.1e-07 PS=9.3e-07
mXI31/XI1/XI41/XI1/MM_instance_280 XI31/XI1/XI41/XI1/NET_009 OP1<3>
+ XI31/XI1/XI41/XI1/NET_010 VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14
+ AS=4.41e-14 PD=9.1e-07 PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_275 VDD! XI31/XI1/NET2 XI31/XI1/XI41/XI1/NET_009
+ VDD! PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06
+ PS=9.1e-07
mXI31/XI1/XI41/XI1/MM_instance_315 XI31/XI1/XI41/S_0<1>
+ XI31/XI1/XI41/XI1/NET_005 VDD! VDD! PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14
+ AS=6.615e-14 PD=1.47e-06 PS=1.54e-06
c_5 C0X<0> 0 0.295485f
c_58 CTRL_BUFF<1> 0 7.10521f
c_178 CTRL_BUFF<0> 0 17.1405f
c_190 OP1<15> 0 2.04018f
c_198 ARITHMETIC_OUT<15> 0 0.632855f
c_212 OP0_TEMP<15> 0 1.36813f
c_216 ALU_PRE_N<15> 0 0.507969f
c_220 CO_N 0 0.611619f
c_226 ALU_PRE<15> 0 0.442976f
c_232 ARITHMETIC_OUT_N<15> 0 0.378835f
c_237 OP1_N<15> 0 0.448871f
c_243 OP0_TEMP_N<15> 0 0.346421f
c_247 V_FLAG 0 0.147533f
c_252 OV1 0 0.353607f
c_256 OV0 0 0.356646f
c_259 C_FLAG 0 0.104743f
c_261 N_FLAG 0 0.236495f
c_266 C0X<2> 0 0.288304f
c_318 CTRL_BUFF<2> 0 7.89399f
c_322 C0X<1> 0 0.352018f
c_512 VSS! 0 39.0184f
c_515 CO 0 0.314304f
c_830 VDD! 0 36.6655f
c_831 CTRL<1> 0 0.193379f
c_833 CTRL<0> 0 0.133232f
c_835 CTRL<2> 0 0.14164f
c_846 OP0<0> 0 0.678849f
c_855 OP1<0> 0 0.917439f
c_858 ALU_OUT<0> 0 0.14958f
c_869 OP0<1> 0 0.676402f
c_879 OP1<1> 0 0.915838f
c_882 ALU_OUT<1> 0 0.149211f
c_893 OP0<2> 0 0.678008f
c_902 OP1<2> 0 1.53063f
c_905 ALU_OUT<2> 0 0.149436f
c_916 OP0<3> 0 0.678177f
c_927 OP1<3> 0 1.52355f
c_930 ALU_OUT<3> 0 0.149281f
c_941 OP0<4> 0 0.676388f
c_950 OP1<4> 0 1.50726f
c_953 ALU_OUT<4> 0 0.149328f
c_964 OP0<5> 0 0.676402f
c_975 OP1<5> 0 1.54135f
c_978 ALU_OUT<5> 0 0.149577f
c_989 OP0<6> 0 0.676421f
c_1000 OP1<6> 0 1.5412f
c_1003 ALU_OUT<6> 0 0.149266f
c_1014 OP0<7> 0 0.676534f
c_1023 OP1<7> 0 1.53052f
c_1026 ALU_OUT<7> 0 0.149577f
c_1037 OP0<8> 0 0.676402f
c_1048 OP1<8> 0 1.54122f
c_1051 ALU_OUT<8> 0 0.149577f
c_1062 OP0<9> 0 0.676402f
c_1073 OP1<9> 0 1.54122f
c_1076 ALU_OUT<9> 0 0.149577f
c_1087 OP0<10> 0 0.676402f
c_1098 OP1<10> 0 1.54126f
c_1101 ALU_OUT<10> 0 0.149174f
c_1112 OP0<11> 0 0.676393f
c_1121 OP1<11> 0 1.53091f
c_1124 ALU_OUT<11> 0 0.149453f
c_1135 OP0<12> 0 0.676503f
c_1146 OP1<12> 0 1.54119f
c_1149 ALU_OUT<12> 0 0.149577f
c_1160 OP0<13> 0 0.676402f
c_1171 OP1<13> 0 1.54122f
c_1174 ALU_OUT<13> 0 0.149577f
c_1185 OP0<14> 0 0.676233f
c_1196 OP1<14> 0 1.54122f
c_1199 ALU_OUT<14> 0 0.149577f
c_1210 OP0<15> 0 0.675337f
c_1214 ALU_OUT<15> 0 0.141273f
c_1221 XI31/XI1/XI40/OP0_TEMP<0> 0 0.608916f
c_1226 XI31/ARITHMETIC_OUT<0> 0 0.422491f
c_1232 XI31/LOGIC_OUT<0> 0 0.540036f
c_1239 XI31/XI1/XI40/OP0_TEMP<1> 0 0.646436f
c_1244 XI31/XI1/XI40/NET16 0 0.544325f
c_1249 XI31/ARITHMETIC_OUT<1> 0 0.432886f
c_1256 XI31/LOGIC_OUT<1> 0 0.491922f
c_1268 XI31/XI1/NET1 0 1.28481f
c_1272 XI31/ARITHMETIC_OUT<2> 0 0.295962f
c_1278 XI31/LOGIC_OUT<2> 0 0.57548f
c_1282 XI31/ARITHMETIC_OUT<3> 0 0.294996f
c_1288 XI31/LOGIC_OUT<3> 0 0.599019f
c_1301 XI31/XI1/NET3 0 1.56755f
c_1305 XI31/ARITHMETIC_OUT<4> 0 0.295381f
c_1311 XI31/LOGIC_OUT<4> 0 0.57159f
c_1315 XI31/ARITHMETIC_OUT<5> 0 0.294125f
c_1321 XI31/LOGIC_OUT<5> 0 0.572979f
c_1325 XI31/ARITHMETIC_OUT<6> 0 0.293232f
c_1331 XI31/LOGIC_OUT<6> 0 0.595831f
c_1346 XI31/XI1/NET12 0 2.08459f
c_1350 XI31/ARITHMETIC_OUT<7> 0 0.294395f
c_1356 XI31/LOGIC_OUT<7> 0 0.586413f
c_1360 XI31/ARITHMETIC_OUT<8> 0 0.294395f
c_1366 XI31/LOGIC_OUT<8> 0 0.586129f
c_1370 XI31/ARITHMETIC_OUT<9> 0 0.294125f
c_1376 XI31/LOGIC_OUT<9> 0 0.586118f
c_1380 XI31/ARITHMETIC_OUT<10> 0 0.293232f
c_1386 XI31/LOGIC_OUT<10> 0 0.595831f
c_1403 XI31/XI1/NET16 0 2.52327f
c_1407 XI31/ARITHMETIC_OUT<11> 0 0.29447f
c_1413 XI31/LOGIC_OUT<11> 0 0.583961f
c_1417 XI31/ARITHMETIC_OUT<12> 0 0.294395f
c_1423 XI31/LOGIC_OUT<12> 0 0.586554f
c_1427 XI31/ARITHMETIC_OUT<13> 0 0.294395f
c_1433 XI31/LOGIC_OUT<13> 0 0.586129f
c_1437 XI31/ARITHMETIC_OUT<14> 0 0.294125f
c_1443 XI31/LOGIC_OUT<14> 0 0.586118f
c_1449 XI31/LOGIC_OUT<15> 0 0.612583f
c_1453 XI31/XI2/ALU_PRE<0> 0 0.297179f
c_1458 XI31/XI2/NET3<15> 0 0.299425f
c_1462 XI31/XI2/ALU_PRE<1> 0 0.297568f
c_1467 XI31/XI2/NET3<14> 0 0.299466f
c_1471 XI31/XI2/ALU_PRE<2> 0 0.295454f
c_1476 XI31/XI2/NET3<13> 0 0.299592f
c_1480 XI31/XI2/ALU_PRE<3> 0 0.296926f
c_1485 XI31/XI2/NET3<12> 0 0.299462f
c_1489 XI31/XI2/ALU_PRE<4> 0 0.295439f
c_1494 XI31/XI2/NET3<11> 0 0.299453f
c_1498 XI31/XI2/ALU_PRE<5> 0 0.295414f
c_1503 XI31/XI2/NET3<10> 0 0.299538f
c_1507 XI31/XI2/ALU_PRE<6> 0 0.297128f
c_1512 XI31/XI2/NET3<9> 0 0.299399f
c_1516 XI31/XI2/ALU_PRE<7> 0 0.295414f
c_1521 XI31/XI2/NET3<8> 0 0.299538f
c_1525 XI31/XI2/ALU_PRE<8> 0 0.295414f
c_1530 XI31/XI2/NET3<7> 0 0.299538f
c_1534 XI31/XI2/ALU_PRE<9> 0 0.295414f
c_1539 XI31/XI2/NET3<6> 0 0.299538f
c_1543 XI31/XI2/ALU_PRE<10> 0 0.297128f
c_1548 XI31/XI2/NET3<5> 0 0.299402f
c_1552 XI31/XI2/ALU_PRE<11> 0 0.295493f
c_1557 XI31/XI2/NET3<4> 0 0.299754f
c_1561 XI31/XI2/ALU_PRE<12> 0 0.295414f
c_1566 XI31/XI2/NET3<3> 0 0.299538f
c_1570 XI31/XI2/ALU_PRE<13> 0 0.295414f
c_1575 XI31/XI2/NET3<2> 0 0.299538f
c_1579 XI31/XI2/ALU_PRE<14> 0 0.295414f
c_1584 XI31/XI2/NET3<1> 0 0.299538f
c_1589 XI31/XI2/NET3<0> 0 0.289882f
c_1593 XI31/XI1/XI40/XI0/NET_001 0 0.373223f
c_1597 XI31/XI1/XI40/XI1/NET_001 0 0.372909f
c_1600 XI31/XI1/XI44/CO_0 0 0.405334f
c_1605 XI31/XI0/XI15/MUX0 0 0.375162f
c_1610 XI31/XI0/XI0/MUX0 0 0.315318f
c_1615 XI31/XI0/XI4/MUX0 0 0.3752f
c_1620 XI31/XI0/XI14/MUX0 0 0.375325f
c_1625 XI31/XI0/XI12/MUX0 0 0.375189f
c_1630 XI31/XI0/XI11/MUX0 0 0.3752f
c_1635 XI31/XI0/XI8/MUX0 0 0.3752f
c_1640 XI31/XI0/XI7/MUX0 0 0.3752f
c_1645 XI31/XI0/XI5/MUX0 0 0.375195f
c_1651 XI31/XI2/XI0<15>/X1 0 0.178886f
c_1655 XI31/XI2/XI0<15>/Z_NEG 0 0.249986f
c_1660 XI31/XI0/XI0/NOR_OUT 0 0.312467f
c_1666 XI31/XI0/XI0/NAND_OUT 0 0.336134f
c_1671 XI31/XI0/XI0/MUX1 0 0.204315f
c_1677 XI31/XI0/XI0/XNOR_OUT 0 0.407702f
c_1680 XI31/XI0/XI0/XI1/NET_000 0 0.241219f
c_1683 XI31/XI0/XI0/XI1/NET_002 0 0.0608951f
c_1688 XI31/XI0/XI0/XI5/Z 0 0.148223f
c_1693 XI31/XI0/XI0/XI4/X1 0 0.200977f
c_1698 XI31/XI0/XI0/XI4/Z_NEG 0 0.16069f
c_1703 XI31/XI0/XI0/XI5/XI0/X1 0 0.175233f
c_1708 XI31/XI0/XI0/XI5/XI0/Z_NEG 0 0.230864f
c_1713 XI31/XI0/XI0/XI3/X1 0 0.282504f
c_1718 XI31/XI0/XI0/XI3/Z_NEG 0 0.213711f
c_1723 XI31/XI2/XI0<14>/X1 0 0.263545f
c_1727 XI31/XI2/XI0<14>/Z_NEG 0 0.232785f
c_1732 XI31/XI0/XI4/NOR_OUT 0 0.312467f
c_1738 XI31/XI0/XI4/NAND_OUT 0 0.336134f
c_1743 XI31/XI0/XI4/MUX1 0 0.204306f
c_1749 XI31/XI0/XI4/XNOR_OUT 0 0.407493f
c_1752 XI31/XI0/XI4/XI1/NET_000 0 0.241219f
c_1755 XI31/XI0/XI4/XI1/NET_002 0 0.0608951f
c_1760 XI31/XI0/XI4/XI5/Z 0 0.148335f
c_1765 XI31/XI0/XI4/XI4/X1 0 0.200962f
c_1770 XI31/XI0/XI4/XI4/Z_NEG 0 0.16061f
c_1775 XI31/XI0/XI4/XI5/XI0/X1 0 0.175287f
c_1780 XI31/XI0/XI4/XI5/XI0/Z_NEG 0 0.23075f
c_1785 XI31/XI0/XI4/XI3/X1 0 0.282504f
c_1790 XI31/XI0/XI4/XI3/Z_NEG 0 0.214063f
c_1795 XI31/XI2/XI0<1>/X1 0 0.263594f
c_1799 XI31/XI2/XI0<1>/Z_NEG 0 0.234698f
c_1804 XI31/XI2/XI0<0>/X1 0 0.266502f
c_1808 XI31/XI2/XI0<0>/Z_NEG 0 0.234698f
c_1813 XI31/XI2/XI0<3>/X1 0 0.26349f
c_1817 XI31/XI2/XI0<3>/Z_NEG 0 0.232765f
c_1822 XI31/XI2/XI0<2>/X1 0 0.263545f
c_1826 XI31/XI2/XI0<2>/Z_NEG 0 0.232765f
c_1831 XI31/XI2/XI0<5>/X1 0 0.263545f
c_1835 XI31/XI2/XI0<5>/Z_NEG 0 0.232785f
c_1840 XI31/XI2/XI0<4>/X1 0 0.263545f
c_1844 XI31/XI2/XI0<4>/Z_NEG 0 0.232785f
c_1849 XI31/XI2/XI0<7>/X1 0 0.263545f
c_1853 XI31/XI2/XI0<7>/Z_NEG 0 0.232785f
c_1858 XI31/XI2/XI0<6>/X1 0 0.263501f
c_1862 XI31/XI2/XI0<6>/Z_NEG 0 0.232785f
c_1867 XI31/XI2/XI0<9>/X1 0 0.263545f
c_1871 XI31/XI2/XI0<9>/Z_NEG 0 0.232785f
c_1876 XI31/XI2/XI0<8>/X1 0 0.263545f
c_1880 XI31/XI2/XI0<8>/Z_NEG 0 0.232785f
c_1885 XI31/XI2/XI0<11>/X1 0 0.263545f
c_1889 XI31/XI2/XI0<11>/Z_NEG 0 0.232785f
c_1894 XI31/XI2/XI0<10>/X1 0 0.263501f
c_1898 XI31/XI2/XI0<10>/Z_NEG 0 0.232785f
c_1903 XI31/XI2/XI0<13>/X1 0 0.263545f
c_1907 XI31/XI2/XI0<13>/Z_NEG 0 0.232785f
c_1912 XI31/XI2/XI0<12>/X1 0 0.263545f
c_1916 XI31/XI2/XI0<12>/Z_NEG 0 0.232785f
c_1921 XI31/XI0/XI16/MUX0 0 0.3752f
c_1926 XI31/XI0/XI15/NOR_OUT 0 0.311639f
c_1932 XI31/XI0/XI15/NAND_OUT 0 0.336898f
c_1937 XI31/XI0/XI15/MUX1 0 0.20779f
c_1943 XI31/XI0/XI15/XNOR_OUT 0 0.407798f
c_1946 XI31/XI0/XI15/XI1/NET_000 0 0.243126f
c_1949 XI31/XI0/XI15/XI1/NET_002 0 0.0609873f
c_1954 XI31/XI0/XI15/XI5/Z 0 0.148335f
c_1959 XI31/XI0/XI15/XI4/X1 0 0.200419f
c_1964 XI31/XI0/XI15/XI4/Z_NEG 0 0.15883f
c_1969 XI31/XI0/XI15/XI5/XI0/X1 0 0.175598f
c_1974 XI31/XI0/XI15/XI5/XI0/Z_NEG 0 0.230656f
c_1979 XI31/XI0/XI15/XI3/X1 0 0.282504f
c_1984 XI31/XI0/XI15/XI3/Z_NEG 0 0.214063f
c_1989 XI31/XI0/XI16/NOR_OUT 0 0.312467f
c_1995 XI31/XI0/XI16/NAND_OUT 0 0.336134f
c_2000 XI31/XI0/XI16/MUX1 0 0.204306f
c_2006 XI31/XI0/XI16/XNOR_OUT 0 0.407493f
c_2009 XI31/XI0/XI16/XI1/NET_000 0 0.241219f
c_2012 XI31/XI0/XI16/XI1/NET_002 0 0.0608951f
c_2017 XI31/XI0/XI16/XI5/Z 0 0.148335f
c_2022 XI31/XI0/XI16/XI4/X1 0 0.200962f
c_2027 XI31/XI0/XI16/XI4/Z_NEG 0 0.16061f
c_2032 XI31/XI0/XI16/XI5/XI0/X1 0 0.175287f
c_2037 XI31/XI0/XI16/XI5/XI0/Z_NEG 0 0.23075f
c_2042 XI31/XI0/XI16/XI3/X1 0 0.282504f
c_2047 XI31/XI0/XI16/XI3/Z_NEG 0 0.214063f
c_2052 XI31/XI0/XI17/MUX0 0 0.375335f
c_2057 XI31/XI0/XI14/NOR_OUT 0 0.313304f
c_2063 XI31/XI0/XI14/NAND_OUT 0 0.336134f
c_2068 XI31/XI0/XI14/MUX1 0 0.207215f
c_2074 XI31/XI0/XI14/XNOR_OUT 0 0.407493f
c_2077 XI31/XI0/XI14/XI1/NET_000 0 0.241219f
c_2080 XI31/XI0/XI14/XI1/NET_002 0 0.0608951f
c_2085 XI31/XI0/XI14/XI5/Z 0 0.148335f
c_2090 XI31/XI0/XI14/XI4/X1 0 0.201032f
c_2095 XI31/XI0/XI14/XI4/Z_NEG 0 0.160478f
c_2100 XI31/XI0/XI14/XI5/XI0/X1 0 0.175254f
c_2105 XI31/XI0/XI14/XI5/XI0/Z_NEG 0 0.230746f
c_2110 XI31/XI0/XI14/XI3/X1 0 0.282504f
c_2115 XI31/XI0/XI14/XI3/Z_NEG 0 0.214063f
c_2120 XI31/XI0/XI17/NOR_OUT 0 0.313304f
c_2126 XI31/XI0/XI17/NAND_OUT 0 0.336134f
c_2131 XI31/XI0/XI17/MUX1 0 0.204338f
c_2137 XI31/XI0/XI17/XNOR_OUT 0 0.407493f
c_2140 XI31/XI0/XI17/XI1/NET_000 0 0.241219f
c_2143 XI31/XI0/XI17/XI1/NET_002 0 0.0608951f
c_2148 XI31/XI0/XI17/XI5/Z 0 0.148335f
c_2153 XI31/XI0/XI17/XI4/X1 0 0.201032f
c_2158 XI31/XI0/XI17/XI4/Z_NEG 0 0.160478f
c_2163 XI31/XI0/XI17/XI5/XI0/X1 0 0.175343f
c_2168 XI31/XI0/XI17/XI5/XI0/Z_NEG 0 0.230746f
c_2173 XI31/XI0/XI17/XI3/X1 0 0.282504f
c_2178 XI31/XI0/XI17/XI3/Z_NEG 0 0.214063f
c_2183 XI31/XI0/XI13/MUX0 0 0.375189f
c_2188 XI31/XI0/XI12/NOR_OUT 0 0.312467f
c_2194 XI31/XI0/XI12/NAND_OUT 0 0.336134f
c_2199 XI31/XI0/XI12/MUX1 0 0.204302f
c_2205 XI31/XI0/XI12/XNOR_OUT 0 0.407493f
c_2208 XI31/XI0/XI12/XI1/NET_000 0 0.241219f
c_2211 XI31/XI0/XI12/XI1/NET_002 0 0.0608951f
c_2216 XI31/XI0/XI12/XI5/Z 0 0.148335f
c_2221 XI31/XI0/XI12/XI4/X1 0 0.200962f
c_2226 XI31/XI0/XI12/XI4/Z_NEG 0 0.16061f
c_2231 XI31/XI0/XI12/XI5/XI0/X1 0 0.175148f
c_2236 XI31/XI0/XI12/XI5/XI0/Z_NEG 0 0.23075f
c_2241 XI31/XI0/XI12/XI3/X1 0 0.282504f
c_2246 XI31/XI0/XI12/XI3/Z_NEG 0 0.214063f
c_2251 XI31/XI0/XI13/NOR_OUT 0 0.312467f
c_2257 XI31/XI0/XI13/NAND_OUT 0 0.336134f
c_2262 XI31/XI0/XI13/MUX1 0 0.204302f
c_2268 XI31/XI0/XI13/XNOR_OUT 0 0.407493f
c_2271 XI31/XI0/XI13/XI1/NET_000 0 0.241219f
c_2274 XI31/XI0/XI13/XI1/NET_002 0 0.0608951f
c_2279 XI31/XI0/XI13/XI5/Z 0 0.148335f
c_2284 XI31/XI0/XI13/XI4/X1 0 0.200962f
c_2289 XI31/XI0/XI13/XI4/Z_NEG 0 0.16061f
c_2294 XI31/XI0/XI13/XI5/XI0/X1 0 0.175148f
c_2299 XI31/XI0/XI13/XI5/XI0/Z_NEG 0 0.23075f
c_2304 XI31/XI0/XI13/XI3/X1 0 0.282504f
c_2309 XI31/XI0/XI13/XI3/Z_NEG 0 0.214063f
c_2314 XI31/XI0/XI18/MUX0 0 0.375195f
c_2319 XI31/XI0/XI11/NOR_OUT 0 0.312467f
c_2325 XI31/XI0/XI11/NAND_OUT 0 0.336134f
c_2330 XI31/XI0/XI11/MUX1 0 0.204306f
c_2336 XI31/XI0/XI11/XNOR_OUT 0 0.407493f
c_2339 XI31/XI0/XI11/XI1/NET_000 0 0.241219f
c_2342 XI31/XI0/XI11/XI1/NET_002 0 0.0608951f
c_2347 XI31/XI0/XI11/XI5/Z 0 0.148335f
c_2352 XI31/XI0/XI11/XI4/X1 0 0.200962f
c_2357 XI31/XI0/XI11/XI4/Z_NEG 0 0.16061f
c_2362 XI31/XI0/XI11/XI5/XI0/X1 0 0.175287f
c_2367 XI31/XI0/XI11/XI5/XI0/Z_NEG 0 0.23075f
c_2372 XI31/XI0/XI11/XI3/X1 0 0.282504f
c_2377 XI31/XI0/XI11/XI3/Z_NEG 0 0.214063f
c_2382 XI31/XI0/XI18/NOR_OUT 0 0.312467f
c_2388 XI31/XI0/XI18/NAND_OUT 0 0.336134f
c_2393 XI31/XI0/XI18/MUX1 0 0.204306f
c_2399 XI31/XI0/XI18/XNOR_OUT 0 0.407493f
c_2402 XI31/XI0/XI18/XI1/NET_000 0 0.241219f
c_2405 XI31/XI0/XI18/XI1/NET_002 0 0.0608951f
c_2410 XI31/XI0/XI18/XI5/Z 0 0.148335f
c_2415 XI31/XI0/XI18/XI4/X1 0 0.200962f
c_2420 XI31/XI0/XI18/XI4/Z_NEG 0 0.16061f
c_2425 XI31/XI0/XI18/XI5/XI0/X1 0 0.175287f
c_2430 XI31/XI0/XI18/XI5/XI0/Z_NEG 0 0.23075f
c_2435 XI31/XI0/XI18/XI3/X1 0 0.282504f
c_2440 XI31/XI0/XI18/XI3/Z_NEG 0 0.214063f
c_2445 XI31/XI0/XI9/MUX0 0 0.3752f
c_2450 XI31/XI0/XI8/NOR_OUT 0 0.312467f
c_2456 XI31/XI0/XI8/NAND_OUT 0 0.336134f
c_2461 XI31/XI0/XI8/MUX1 0 0.204306f
c_2467 XI31/XI0/XI8/XNOR_OUT 0 0.407493f
c_2470 XI31/XI0/XI8/XI1/NET_000 0 0.241219f
c_2473 XI31/XI0/XI8/XI1/NET_002 0 0.0608951f
c_2478 XI31/XI0/XI8/XI5/Z 0 0.148335f
c_2483 XI31/XI0/XI8/XI4/X1 0 0.200962f
c_2488 XI31/XI0/XI8/XI4/Z_NEG 0 0.16061f
c_2493 XI31/XI0/XI8/XI5/XI0/X1 0 0.175287f
c_2498 XI31/XI0/XI8/XI5/XI0/Z_NEG 0 0.23075f
c_2503 XI31/XI0/XI8/XI3/X1 0 0.282504f
c_2508 XI31/XI0/XI8/XI3/Z_NEG 0 0.214063f
c_2513 XI31/XI0/XI9/NOR_OUT 0 0.312467f
c_2519 XI31/XI0/XI9/NAND_OUT 0 0.336134f
c_2524 XI31/XI0/XI9/MUX1 0 0.204306f
c_2530 XI31/XI0/XI9/XNOR_OUT 0 0.407493f
c_2533 XI31/XI0/XI9/XI1/NET_000 0 0.241219f
c_2536 XI31/XI0/XI9/XI1/NET_002 0 0.0608951f
c_2541 XI31/XI0/XI9/XI5/Z 0 0.148335f
c_2546 XI31/XI0/XI9/XI4/X1 0 0.200962f
c_2551 XI31/XI0/XI9/XI4/Z_NEG 0 0.16061f
c_2556 XI31/XI0/XI9/XI5/XI0/X1 0 0.175287f
c_2561 XI31/XI0/XI9/XI5/XI0/Z_NEG 0 0.23075f
c_2566 XI31/XI0/XI9/XI3/X1 0 0.282504f
c_2571 XI31/XI0/XI9/XI3/Z_NEG 0 0.214063f
c_2576 XI31/XI0/XI10/MUX0 0 0.375171f
c_2581 XI31/XI0/XI7/NOR_OUT 0 0.312467f
c_2587 XI31/XI0/XI7/NAND_OUT 0 0.336134f
c_2592 XI31/XI0/XI7/MUX1 0 0.204306f
c_2598 XI31/XI0/XI7/XNOR_OUT 0 0.407493f
c_2601 XI31/XI0/XI7/XI1/NET_000 0 0.241219f
c_2604 XI31/XI0/XI7/XI1/NET_002 0 0.0608951f
c_2609 XI31/XI0/XI7/XI5/Z 0 0.148335f
c_2614 XI31/XI0/XI7/XI4/X1 0 0.200962f
c_2619 XI31/XI0/XI7/XI4/Z_NEG 0 0.16061f
c_2624 XI31/XI0/XI7/XI5/XI0/X1 0 0.175287f
c_2629 XI31/XI0/XI7/XI5/XI0/Z_NEG 0 0.23075f
c_2634 XI31/XI0/XI7/XI3/X1 0 0.282504f
c_2639 XI31/XI0/XI7/XI3/Z_NEG 0 0.214063f
c_2644 XI31/XI0/XI10/NOR_OUT 0 0.312467f
c_2650 XI31/XI0/XI10/NAND_OUT 0 0.336134f
c_2655 XI31/XI0/XI10/MUX1 0 0.204306f
c_2661 XI31/XI0/XI10/XNOR_OUT 0 0.407493f
c_2664 XI31/XI0/XI10/XI1/NET_000 0 0.241219f
c_2667 XI31/XI0/XI10/XI1/NET_002 0 0.0608951f
c_2672 XI31/XI0/XI10/XI5/Z 0 0.148335f
c_2677 XI31/XI0/XI10/XI4/X1 0 0.200962f
c_2682 XI31/XI0/XI10/XI4/Z_NEG 0 0.16061f
c_2687 XI31/XI0/XI10/XI5/XI0/X1 0 0.175077f
c_2692 XI31/XI0/XI10/XI5/XI0/Z_NEG 0 0.23075f
c_2697 XI31/XI0/XI10/XI3/X1 0 0.282504f
c_2702 XI31/XI0/XI10/XI3/Z_NEG 0 0.214063f
c_2707 XI31/XI0/XI6/MUX0 0 0.3752f
c_2712 XI31/XI0/XI5/NOR_OUT 0 0.312467f
c_2718 XI31/XI0/XI5/NAND_OUT 0 0.336134f
c_2723 XI31/XI0/XI5/MUX1 0 0.204306f
c_2729 XI31/XI0/XI5/XNOR_OUT 0 0.407493f
c_2732 XI31/XI0/XI5/XI1/NET_000 0 0.241219f
c_2735 XI31/XI0/XI5/XI1/NET_002 0 0.0608951f
c_2740 XI31/XI0/XI5/XI5/Z 0 0.148335f
c_2745 XI31/XI0/XI5/XI4/X1 0 0.200962f
c_2750 XI31/XI0/XI5/XI4/Z_NEG 0 0.16061f
c_2755 XI31/XI0/XI5/XI5/XI0/X1 0 0.175287f
c_2760 XI31/XI0/XI5/XI5/XI0/Z_NEG 0 0.23075f
c_2765 XI31/XI0/XI5/XI3/X1 0 0.282504f
c_2770 XI31/XI0/XI5/XI3/Z_NEG 0 0.214063f
c_2775 XI31/XI0/XI6/NOR_OUT 0 0.312467f
c_2781 XI31/XI0/XI6/NAND_OUT 0 0.336134f
c_2786 XI31/XI0/XI6/MUX1 0 0.204306f
c_2792 XI31/XI0/XI6/XNOR_OUT 0 0.407493f
c_2795 XI31/XI0/XI6/XI1/NET_000 0 0.241219f
c_2798 XI31/XI0/XI6/XI1/NET_002 0 0.0608951f
c_2803 XI31/XI0/XI6/XI5/Z 0 0.148335f
c_2808 XI31/XI0/XI6/XI4/X1 0 0.200962f
c_2813 XI31/XI0/XI6/XI4/Z_NEG 0 0.16061f
c_2818 XI31/XI0/XI6/XI5/XI0/X1 0 0.175287f
c_2823 XI31/XI0/XI6/XI5/XI0/Z_NEG 0 0.23075f
c_2828 XI31/XI0/XI6/XI3/X1 0 0.282504f
c_2833 XI31/XI0/XI6/XI3/Z_NEG 0 0.214063f
c_2835 XI31/XI1/XI40/XI9/NET_000 0 0.243584f
c_2837 XI31/XI1/XI40/XI9/NET_003 0 0.0932618f
c_2839 XI31/XI1/XI40/XI10/NET_000 0 0.226373f
c_2841 XI31/XI1/XI40/XI10/NET_003 0 0.0936387f
c_2842 XI31/XI1/XI40/XI0/NET_002 0 0.163564f
c_2844 XI31/XI1/XI40/XI0/NET_008 0 0.137733f
c_2845 XI31/XI1/XI40/XI0/NET_006 0 0.150238f
c_2847 XI31/XI1/XI40/XI0/NET_011 0 0.137533f
c_2850 XI31/XI1/XI40/XI0/NET_005 0 0.314105f
c_2851 XI31/XI1/XI40/XI1/NET_002 0 0.166092f
c_2853 XI31/XI1/XI40/XI1/NET_008 0 0.137733f
c_2854 XI31/XI1/XI40/XI1/NET_006 0 0.124964f
c_2856 XI31/XI1/XI40/XI1/NET_011 0 0.137653f
c_2859 XI31/XI1/XI40/XI1/NET_005 0 0.328321f
c_2869 XI31/XI1/XI44/OP0_TEMP<0> 0 0.954291f
c_2873 XI31/XI1/XI44/S_0<0> 0 0.370804f
c_2877 XI31/XI1/XI44/S_1<0> 0 0.398806f
c_2888 XI31/XI1/XI44/OP0_TEMP<1> 0 1.04528f
c_2893 XI31/XI1/XI44/NET16 0 0.540852f
c_2898 XI31/XI1/XI44/NET36 0 0.575741f
c_2902 XI31/XI1/XI44/S_0<1> 0 0.400002f
c_2906 XI31/XI1/XI44/S_1<1> 0 0.395896f
c_2917 XI31/XI1/XI44/OP0_TEMP<2> 0 1.04522f
c_2922 XI31/XI1/XI44/NET21 0 0.541791f
c_2927 XI31/XI1/XI44/NET41 0 0.578145f
c_2931 XI31/XI1/XI44/S_0<2> 0 0.397608f
c_2935 XI31/XI1/XI44/S_1<2> 0 0.395869f
c_2946 XI31/XI1/XI44/OP0_TEMP<3> 0 1.04522f
c_2951 XI31/XI1/XI44/NET26 0 0.541614f
c_2956 XI31/XI1/XI44/NET46 0 0.57979f
c_2960 XI31/XI1/XI44/S_0<3> 0 0.396087f
c_2964 XI31/XI1/XI44/S_1<3> 0 0.395216f
c_2969 XI31/XI1/XI44/NET2 0 0.534484f
c_2974 XI31/XI1/XI44/NET1 0 0.578432f
c_2978 XI31/XI1/XI44/S_0<4> 0 0.397783f
c_2982 XI31/XI1/XI44/S_1<4> 0 0.367152f
c_2986 XI31/XI1/XI44/CO_1 0 0.301887f
c_2989 XI31/XI1/XI44/XI32/NET_001 0 0.452352f
c_2993 XI31/XI1/XI44/XI5/NET_001 0 0.344941f
c_2997 XI31/XI1/XI44/XI0/NET_001 0 0.342417f
c_3001 XI31/XI1/XI44/XI6/NET_001 0 0.374788f
c_3005 XI31/XI1/XI44/XI1/NET_001 0 0.375633f
c_3009 XI31/XI1/XI44/XI7/NET_001 0 0.374748f
c_3013 XI31/XI1/XI44/XI2/NET_001 0 0.375633f
c_3017 XI31/XI1/XI44/XI8/NET_001 0 0.374748f
c_3021 XI31/XI1/XI44/XI3/NET_001 0 0.375633f
c_3025 XI31/XI1/XI44/XI33/NET_001 0 0.379841f
c_3030 XI31/XI1/XI44/XI17/X1 0 0.16862f
c_3034 XI31/XI1/XI44/XI17/Z_NEG 0 0.234387f
c_3039 XI31/XI1/XI44/XI25/X1 0 0.166163f
c_3043 XI31/XI1/XI44/XI25/Z_NEG 0 0.23521f
c_3048 XI31/XI1/XI44/XI26/X1 0 0.166248f
c_3052 XI31/XI1/XI44/XI26/Z_NEG 0 0.23521f
c_3057 XI31/XI1/XI44/XI24/X1 0 0.166098f
c_3061 XI31/XI1/XI44/XI24/Z_NEG 0 0.23492f
c_3066 XI31/XI1/XI44/XI35/X1 0 0.166248f
c_3070 XI31/XI1/XI44/XI35/Z_NEG 0 0.235128f
c_3073 XI31/XI1/XI44/XI18/X1 0 0.327698f
c_3077 XI31/XI1/XI44/XI18/Z_NEG 0 0.233263f
c_3079 XI31/XI1/XI44/XI9/NET_000 0 0.227217f
c_3081 XI31/XI1/XI44/XI9/NET_003 0 0.0936829f
c_3083 XI31/XI1/XI44/XI10/NET_000 0 0.226354f
c_3085 XI31/XI1/XI44/XI10/NET_003 0 0.0934226f
c_3087 XI31/XI1/XI44/XI11/NET_000 0 0.226373f
c_3089 XI31/XI1/XI44/XI11/NET_003 0 0.0936387f
c_3091 XI31/XI1/XI44/XI12/NET_000 0 0.226871f
c_3093 XI31/XI1/XI44/XI12/NET_003 0 0.0939347f
c_3095 XI31/XI1/XI44/XI34/NET_000 0 0.232446f
c_3097 XI31/XI1/XI44/XI34/NET_003 0 0.0946896f
c_3098 XI31/XI1/XI44/XI5/NET_002 0 0.160314f
c_3100 XI31/XI1/XI44/XI5/NET_008 0 0.135348f
c_3102 XI31/XI1/XI44/XI5/NET_006 0 0.195256f
c_3105 XI31/XI1/XI44/XI5/NET_011 0 0.0325446f
c_3109 XI31/XI1/XI44/XI5/NET_005 0 0.334433f
c_3111 XI31/XI1/XI44/XI0/NET_002 0 0.0551793f
c_3112 XI31/XI1/XI44/XI0/NET_008 0 0.230781f
c_3113 XI31/XI1/XI44/XI0/NET_006 0 0.1575f
c_3115 XI31/XI1/XI44/XI0/NET_011 0 0.135307f
c_3118 XI31/XI1/XI44/XI0/NET_005 0 0.309048f
c_3119 XI31/XI1/XI44/XI6/NET_002 0 0.160314f
c_3120 XI31/XI1/XI44/XI6/NET_008 0 0.230799f
c_3122 XI31/XI1/XI44/XI6/NET_006 0 0.195203f
c_3124 XI31/XI1/XI44/XI6/NET_011 0 0.135422f
c_3128 XI31/XI1/XI44/XI6/NET_005 0 0.336229f
c_3129 XI31/XI1/XI44/XI1/NET_002 0 0.164577f
c_3130 XI31/XI1/XI44/XI1/NET_008 0 0.230781f
c_3131 XI31/XI1/XI44/XI1/NET_006 0 0.131676f
c_3133 XI31/XI1/XI44/XI1/NET_011 0 0.135474f
c_3136 XI31/XI1/XI44/XI1/NET_005 0 0.323429f
c_3137 XI31/XI1/XI44/XI7/NET_002 0 0.160314f
c_3138 XI31/XI1/XI44/XI7/NET_008 0 0.230799f
c_3140 XI31/XI1/XI44/XI7/NET_006 0 0.195203f
c_3142 XI31/XI1/XI44/XI7/NET_011 0 0.135422f
c_3146 XI31/XI1/XI44/XI7/NET_005 0 0.336047f
c_3147 XI31/XI1/XI44/XI2/NET_002 0 0.164855f
c_3148 XI31/XI1/XI44/XI2/NET_008 0 0.230781f
c_3149 XI31/XI1/XI44/XI2/NET_006 0 0.131676f
c_3151 XI31/XI1/XI44/XI2/NET_011 0 0.135474f
c_3154 XI31/XI1/XI44/XI2/NET_005 0 0.323429f
c_3155 XI31/XI1/XI44/XI8/NET_002 0 0.160314f
c_3156 XI31/XI1/XI44/XI8/NET_008 0 0.230799f
c_3158 XI31/XI1/XI44/XI8/NET_006 0 0.195203f
c_3160 XI31/XI1/XI44/XI8/NET_011 0 0.135422f
c_3164 XI31/XI1/XI44/XI8/NET_005 0 0.336047f
c_3165 XI31/XI1/XI44/XI3/NET_002 0 0.164855f
c_3166 XI31/XI1/XI44/XI3/NET_008 0 0.230781f
c_3167 XI31/XI1/XI44/XI3/NET_006 0 0.131676f
c_3169 XI31/XI1/XI44/XI3/NET_011 0 0.135474f
c_3172 XI31/XI1/XI44/XI3/NET_005 0 0.323429f
c_3173 XI31/XI1/XI44/XI32/NET_002 0 0.160598f
c_3174 XI31/XI1/XI44/XI32/NET_008 0 0.230781f
c_3176 XI31/XI1/XI44/XI32/NET_006 0 0.195785f
c_3178 XI31/XI1/XI44/XI32/NET_011 0 0.135422f
c_3182 XI31/XI1/XI44/XI32/NET_005 0 0.336047f
c_3183 XI31/XI1/XI44/XI33/NET_002 0 0.213117f
c_3184 XI31/XI1/XI44/XI33/NET_008 0 0.230566f
c_3186 XI31/XI1/XI44/XI33/NET_006 0 0.0864539f
c_3188 XI31/XI1/XI44/XI33/NET_011 0 0.135368f
c_3191 XI31/XI1/XI44/XI33/NET_005 0 0.322144f
c_3201 XI31/XI1/XI43/OP0_TEMP<0> 0 0.9543f
c_3205 XI31/XI1/XI43/S_0<0> 0 0.372927f
c_3209 XI31/XI1/XI43/S_1<0> 0 0.397683f
c_3220 XI31/XI1/XI43/OP0_TEMP<1> 0 1.04522f
c_3225 XI31/XI1/XI43/NET16 0 0.541791f
c_3230 XI31/XI1/XI43/NET36 0 0.578145f
c_3234 XI31/XI1/XI43/S_0<1> 0 0.397608f
c_3238 XI31/XI1/XI43/S_1<1> 0 0.395869f
c_3249 XI31/XI1/XI43/OP0_TEMP<2> 0 1.04522f
c_3254 XI31/XI1/XI43/NET21 0 0.541791f
c_3259 XI31/XI1/XI43/NET41 0 0.57979f
c_3263 XI31/XI1/XI43/S_0<2> 0 0.396087f
c_3267 XI31/XI1/XI43/S_1<2> 0 0.395216f
c_3278 XI31/XI1/NET18 0 1.04213f
c_3283 XI31/XI1/XI43/NET26 0 0.541791f
c_3288 XI31/XI1/XI43/NET46 0 0.578432f
c_3292 XI31/XI1/XI43/S_0<3> 0 0.397608f
c_3296 XI31/XI1/XI43/S_1<3> 0 0.367115f
c_3299 XI31/XI1/XI43/CO_0 0 0.378317f
c_3303 XI31/XI1/XI43/CO_1 0 0.287569f
c_3306 XI31/XI1/XI43/XI8/NET_001 0 0.452352f
c_3310 XI31/XI1/XI43/XI5/NET_001 0 0.344929f
c_3314 XI31/XI1/XI43/XI0/NET_001 0 0.342523f
c_3318 XI31/XI1/XI43/XI6/NET_001 0 0.374748f
c_3322 XI31/XI1/XI43/XI1/NET_001 0 0.375633f
c_3326 XI31/XI1/XI43/XI7/NET_001 0 0.374748f
c_3330 XI31/XI1/XI43/XI2/NET_001 0 0.375633f
c_3334 XI31/XI1/XI43/XI3/NET_001 0 0.375554f
c_3339 XI31/XI1/XI43/XI17/X1 0 0.166127f
c_3343 XI31/XI1/XI43/XI17/Z_NEG 0 0.23521f
c_3348 XI31/XI1/XI43/XI25/X1 0 0.166248f
c_3352 XI31/XI1/XI43/XI25/Z_NEG 0 0.23521f
c_3357 XI31/XI1/XI43/XI26/X1 0 0.166098f
c_3361 XI31/XI1/XI43/XI26/Z_NEG 0 0.23492f
c_3366 XI31/XI1/XI43/XI24/X1 0 0.166248f
c_3370 XI31/XI1/XI43/XI24/Z_NEG 0 0.234788f
c_3373 XI31/XI1/XI43/XI18/X1 0 0.317402f
c_3376 XI31/XI1/XI43/XI18/Z_NEG 0 0.29038f
c_3378 XI31/XI1/XI43/XI9/NET_000 0 0.227084f
c_3380 XI31/XI1/XI43/XI9/NET_003 0 0.0932152f
c_3382 XI31/XI1/XI43/XI10/NET_000 0 0.226373f
c_3384 XI31/XI1/XI43/XI10/NET_003 0 0.0936387f
c_3386 XI31/XI1/XI43/XI11/NET_000 0 0.226398f
c_3388 XI31/XI1/XI43/XI11/NET_003 0 0.0936387f
c_3390 XI31/XI1/XI43/XI12/NET_000 0 0.226398f
c_3392 XI31/XI1/XI43/XI12/NET_003 0 0.0936387f
c_3393 XI31/XI1/XI43/XI5/NET_002 0 0.160314f
c_3395 XI31/XI1/XI43/XI5/NET_008 0 0.135348f
c_3397 XI31/XI1/XI43/XI5/NET_006 0 0.195256f
c_3400 XI31/XI1/XI43/XI5/NET_011 0 0.0325446f
c_3404 XI31/XI1/XI43/XI5/NET_005 0 0.330897f
c_3406 XI31/XI1/XI43/XI0/NET_002 0 0.0551793f
c_3407 XI31/XI1/XI43/XI0/NET_008 0 0.230781f
c_3408 XI31/XI1/XI43/XI0/NET_006 0 0.1575f
c_3410 XI31/XI1/XI43/XI0/NET_011 0 0.135307f
c_3413 XI31/XI1/XI43/XI0/NET_005 0 0.311586f
c_3414 XI31/XI1/XI43/XI6/NET_002 0 0.160314f
c_3415 XI31/XI1/XI43/XI6/NET_008 0 0.230799f
c_3417 XI31/XI1/XI43/XI6/NET_006 0 0.195203f
c_3419 XI31/XI1/XI43/XI6/NET_011 0 0.135422f
c_3423 XI31/XI1/XI43/XI6/NET_005 0 0.336047f
c_3424 XI31/XI1/XI43/XI1/NET_002 0 0.164855f
c_3425 XI31/XI1/XI43/XI1/NET_008 0 0.230781f
c_3426 XI31/XI1/XI43/XI1/NET_006 0 0.131676f
c_3428 XI31/XI1/XI43/XI1/NET_011 0 0.135474f
c_3431 XI31/XI1/XI43/XI1/NET_005 0 0.323429f
c_3432 XI31/XI1/XI43/XI7/NET_002 0 0.160314f
c_3433 XI31/XI1/XI43/XI7/NET_008 0 0.230799f
c_3435 XI31/XI1/XI43/XI7/NET_006 0 0.195203f
c_3437 XI31/XI1/XI43/XI7/NET_011 0 0.135422f
c_3441 XI31/XI1/XI43/XI7/NET_005 0 0.336047f
c_3442 XI31/XI1/XI43/XI2/NET_002 0 0.164855f
c_3443 XI31/XI1/XI43/XI2/NET_008 0 0.230781f
c_3444 XI31/XI1/XI43/XI2/NET_006 0 0.131676f
c_3446 XI31/XI1/XI43/XI2/NET_011 0 0.135474f
c_3449 XI31/XI1/XI43/XI2/NET_005 0 0.323429f
c_3450 XI31/XI1/XI43/XI8/NET_002 0 0.160598f
c_3451 XI31/XI1/XI43/XI8/NET_008 0 0.230781f
c_3453 XI31/XI1/XI43/XI8/NET_006 0 0.195785f
c_3455 XI31/XI1/XI43/XI8/NET_011 0 0.135422f
c_3459 XI31/XI1/XI43/XI8/NET_005 0 0.336047f
c_3460 XI31/XI1/XI43/XI3/NET_002 0 0.164855f
c_3461 XI31/XI1/XI43/XI3/NET_008 0 0.230781f
c_3462 XI31/XI1/XI43/XI3/NET_006 0 0.131676f
c_3464 XI31/XI1/XI43/XI3/NET_011 0 0.135474f
c_3467 XI31/XI1/XI43/XI3/NET_005 0 0.323429f
c_3477 XI31/XI1/XI42/OP0_TEMP<0> 0 0.956885f
c_3481 XI31/XI1/XI42/S_0<0> 0 0.37106f
c_3485 XI31/XI1/XI42/S_1<0> 0 0.395903f
c_3496 XI31/XI1/XI42/OP0_TEMP<1> 0 1.04523f
c_3501 XI31/XI1/XI42/NET16 0 0.541399f
c_3506 XI31/XI1/XI42/NET36 0 0.579164f
c_3510 XI31/XI1/XI42/S_0<1> 0 0.396212f
c_3514 XI31/XI1/XI42/S_1<1> 0 0.395216f
c_3525 XI31/XI1/NET11 0 1.04213f
c_3530 XI31/XI1/XI42/NET21 0 0.542313f
c_3535 XI31/XI1/XI42/NET41 0 0.578432f
c_3539 XI31/XI1/XI42/S_0<2> 0 0.397608f
c_3543 XI31/XI1/XI42/S_1<2> 0 0.367115f
c_3546 XI31/XI1/XI42/CO_0 0 0.378317f
c_3550 XI31/XI1/XI42/CO_1 0 0.287569f
c_3553 XI31/XI1/XI42/XI7/NET_001 0 0.452352f
c_3557 XI31/XI1/XI42/XI5/NET_001 0 0.344386f
c_3561 XI31/XI1/XI42/XI0/NET_001 0 0.34234f
c_3565 XI31/XI1/XI42/XI6/NET_001 0 0.374748f
c_3569 XI31/XI1/XI42/XI1/NET_001 0 0.375633f
c_3573 XI31/XI1/XI42/XI2/NET_001 0 0.375554f
c_3578 XI31/XI1/XI42/XI17/X1 0 0.166127f
c_3582 XI31/XI1/XI42/XI17/Z_NEG 0 0.23521f
c_3587 XI31/XI1/XI42/XI25/X1 0 0.166098f
c_3591 XI31/XI1/XI42/XI25/Z_NEG 0 0.23492f
c_3596 XI31/XI1/XI42/XI26/X1 0 0.166248f
c_3600 XI31/XI1/XI42/XI26/Z_NEG 0 0.234788f
c_3603 XI31/XI1/XI42/XI18/X1 0 0.317402f
c_3606 XI31/XI1/XI42/XI18/Z_NEG 0 0.290383f
c_3608 XI31/XI1/XI42/XI9/NET_000 0 0.231392f
c_3610 XI31/XI1/XI42/XI9/NET_003 0 0.0937109f
c_3612 XI31/XI1/XI42/XI10/NET_000 0 0.230266f
c_3614 XI31/XI1/XI42/XI10/NET_003 0 0.0936387f
c_3616 XI31/XI1/XI42/XI11/NET_000 0 0.226407f
c_3618 XI31/XI1/XI42/XI11/NET_003 0 0.093535f
c_3619 XI31/XI1/XI42/XI5/NET_002 0 0.160323f
c_3621 XI31/XI1/XI42/XI5/NET_008 0 0.135348f
c_3623 XI31/XI1/XI42/XI5/NET_006 0 0.18649f
c_3626 XI31/XI1/XI42/XI5/NET_011 0 0.0322267f
c_3630 XI31/XI1/XI42/XI5/NET_005 0 0.322441f
c_3632 XI31/XI1/XI42/XI0/NET_002 0 0.0532369f
c_3633 XI31/XI1/XI42/XI0/NET_008 0 0.230781f
c_3634 XI31/XI1/XI42/XI0/NET_006 0 0.162998f
c_3636 XI31/XI1/XI42/XI0/NET_011 0 0.135336f
c_3639 XI31/XI1/XI42/XI0/NET_005 0 0.307665f
c_3640 XI31/XI1/XI42/XI6/NET_002 0 0.160314f
c_3641 XI31/XI1/XI42/XI6/NET_008 0 0.230799f
c_3643 XI31/XI1/XI42/XI6/NET_006 0 0.195203f
c_3645 XI31/XI1/XI42/XI6/NET_011 0 0.135422f
c_3649 XI31/XI1/XI42/XI6/NET_005 0 0.336047f
c_3650 XI31/XI1/XI42/XI1/NET_002 0 0.162547f
c_3651 XI31/XI1/XI42/XI1/NET_008 0 0.230781f
c_3652 XI31/XI1/XI42/XI1/NET_006 0 0.131676f
c_3654 XI31/XI1/XI42/XI1/NET_011 0 0.135474f
c_3657 XI31/XI1/XI42/XI1/NET_005 0 0.323429f
c_3658 XI31/XI1/XI42/XI7/NET_002 0 0.160598f
c_3659 XI31/XI1/XI42/XI7/NET_008 0 0.230781f
c_3661 XI31/XI1/XI42/XI7/NET_006 0 0.195785f
c_3663 XI31/XI1/XI42/XI7/NET_011 0 0.135422f
c_3667 XI31/XI1/XI42/XI7/NET_005 0 0.336047f
c_3668 XI31/XI1/XI42/XI2/NET_002 0 0.164855f
c_3669 XI31/XI1/XI42/XI2/NET_008 0 0.230781f
c_3670 XI31/XI1/XI42/XI2/NET_006 0 0.131676f
c_3672 XI31/XI1/XI42/XI2/NET_011 0 0.135474f
c_3675 XI31/XI1/XI42/XI2/NET_005 0 0.323429f
c_3685 XI31/XI1/XI41/OP0_TEMP<0> 0 0.956732f
c_3689 XI31/XI1/XI41/S_0<0> 0 0.368921f
c_3693 XI31/XI1/XI41/S_1<0> 0 0.388667f
c_3704 XI31/XI1/NET2 0 1.04214f
c_3709 XI31/XI1/XI41/NET16 0 0.541791f
c_3714 XI31/XI1/XI41/NET36 0 0.578529f
c_3718 XI31/XI1/XI41/S_0<1> 0 0.397592f
c_3722 XI31/XI1/XI41/S_1<1> 0 0.366498f
c_3725 XI31/XI1/XI41/CO_0 0 0.378323f
c_3729 XI31/XI1/XI41/CO_1 0 0.287596f
c_3732 XI31/XI1/XI41/XI6/NET_001 0 0.452187f
c_3736 XI31/XI1/XI41/XI5/NET_001 0 0.344553f
c_3740 XI31/XI1/XI41/XI0/NET_001 0 0.342469f
c_3744 XI31/XI1/XI41/XI1/NET_001 0 0.375554f
c_3749 XI31/XI1/XI41/XI17/X1 0 0.166392f
c_3753 XI31/XI1/XI41/XI17/Z_NEG 0 0.236592f
c_3758 XI31/XI1/XI41/XI25/X1 0 0.166627f
c_3762 XI31/XI1/XI41/XI25/Z_NEG 0 0.236332f
c_3765 XI31/XI1/XI41/XI18/X1 0 0.317402f
c_3768 XI31/XI1/XI41/XI18/Z_NEG 0 0.290362f
c_3770 XI31/XI1/XI41/XI9/NET_000 0 0.233834f
c_3772 XI31/XI1/XI41/XI9/NET_003 0 0.0945206f
c_3774 XI31/XI1/XI41/XI10/NET_000 0 0.226725f
c_3776 XI31/XI1/XI41/XI10/NET_003 0 0.0940656f
c_3777 XI31/XI1/XI41/XI5/NET_002 0 0.160314f
c_3779 XI31/XI1/XI41/XI5/NET_008 0 0.135348f
c_3781 XI31/XI1/XI41/XI5/NET_006 0 0.195251f
c_3784 XI31/XI1/XI41/XI5/NET_011 0 0.0322267f
c_3788 XI31/XI1/XI41/XI5/NET_005 0 0.330887f
c_3790 XI31/XI1/XI41/XI0/NET_002 0 0.0546364f
c_3791 XI31/XI1/XI41/XI0/NET_008 0 0.230781f
c_3792 XI31/XI1/XI41/XI0/NET_006 0 0.163506f
c_3794 XI31/XI1/XI41/XI0/NET_011 0 0.135336f
c_3797 XI31/XI1/XI41/XI0/NET_005 0 0.308116f
c_3798 XI31/XI1/XI41/XI6/NET_002 0 0.160429f
c_3799 XI31/XI1/XI41/XI6/NET_008 0 0.230781f
c_3801 XI31/XI1/XI41/XI6/NET_006 0 0.185513f
c_3803 XI31/XI1/XI41/XI6/NET_011 0 0.135422f
c_3807 XI31/XI1/XI41/XI6/NET_005 0 0.327506f
c_3808 XI31/XI1/XI41/XI1/NET_002 0 0.164855f
c_3809 XI31/XI1/XI41/XI1/NET_008 0 0.230781f
c_3810 XI31/XI1/XI41/XI1/NET_006 0 0.131676f
c_3812 XI31/XI1/XI41/XI1/NET_011 0 0.135474f
c_3815 XI31/XI1/XI41/XI1/NET_005 0 0.323429f
*
.include "./ALU.pex.netlist.ALU.pxi"
*
.ends
*
*
