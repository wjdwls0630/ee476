.GLOBAL vdd! vss!


.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2

* File: LFSR.pex.netlist
* Created: Tue Nov  9 02:22:27 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.subckt LFSR  RST CLK STATE<0> STATE<1> STATE<2> STATE<3> STATE<4>
+ STATE<5> STATE<6> STATE<7> STATE<8> STATE<9> STATE<10> STATE<11> STATE<12>
+ STATE<13> STATE<14> STATE<15>
* 
mXxor0.XI0.XI2.MNMOS0 XXOR0.XI0.XI2.NET2 XXOR0.XI0.NET2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI2.MNMOS1 XXOR0.NET1 XXOR0.XI0.NET3 XXOR0.XI0.XI2.NET2 VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI0.XI2.MPMOS0 XXOR0.NET1 XXOR0.XI0.NET2 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI2.MPMOS1 XXOR0.NET1 XXOR0.XI0.NET3 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI0.MNMOS0 XXOR0.XI0.XI0.NET2 STATE<3> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI0.MNMOS1 XXOR0.XI0.NET2 XXOR0.XI0.NET1 XXOR0.XI0.XI0.NET2 VSS!
+ NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI0.XI0.MPMOS0 XXOR0.XI0.NET2 STATE<3> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI0.MPMOS1 XXOR0.XI0.NET2 XXOR0.XI0.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.Xnand0.MNMOS0 XXOR0.XI0.XNAND0.NET2 STATE<3> VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.Xnand0.MNMOS1 XXOR0.XI0.NET1 STATE<5> XXOR0.XI0.XNAND0.NET2 VSS!
+ NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI0.Xnand0.MPMOS0 XXOR0.XI0.NET1 STATE<3> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.Xnand0.MPMOS1 XXOR0.XI0.NET1 STATE<5> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI1.MNMOS0 XXOR0.XI0.XI1.NET2 XXOR0.XI0.NET1 VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI1.MNMOS1 XXOR0.XI0.NET3 STATE<5> XXOR0.XI0.XI1.NET2 VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI0.XI1.MPMOS0 XXOR0.XI0.NET3 XXOR0.XI0.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI0.XI1.MPMOS1 XXOR0.XI0.NET3 STATE<5> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI2.MNMOS0 XXOR0.XI1.XI2.NET2 XXOR0.XI1.NET2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI2.MNMOS1 XXOR0.NET2 XXOR0.XI1.NET3 XXOR0.XI1.XI2.NET2 VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI1.XI2.MPMOS0 XXOR0.NET2 XXOR0.XI1.NET2 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI2.MPMOS1 XXOR0.NET2 XXOR0.XI1.NET3 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI0.MNMOS0 XXOR0.XI1.XI0.NET2 STATE<2> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI0.MNMOS1 XXOR0.XI1.NET2 XXOR0.XI1.NET1 XXOR0.XI1.XI0.NET2 VSS!
+ NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI1.XI0.MPMOS0 XXOR0.XI1.NET2 STATE<2> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI0.MPMOS1 XXOR0.XI1.NET2 XXOR0.XI1.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.Xnand0.MNMOS0 XXOR0.XI1.XNAND0.NET2 STATE<2> VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.Xnand0.MNMOS1 XXOR0.XI1.NET1 XXOR0.NET1 XXOR0.XI1.XNAND0.NET2 VSS!
+ NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI1.Xnand0.MPMOS0 XXOR0.XI1.NET1 STATE<2> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.Xnand0.MPMOS1 XXOR0.XI1.NET1 XXOR0.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI1.MNMOS0 XXOR0.XI1.XI1.NET2 XXOR0.XI1.NET1 VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI1.MNMOS1 XXOR0.XI1.NET3 XXOR0.NET1 XXOR0.XI1.XI1.NET2 VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI1.XI1.MPMOS0 XXOR0.XI1.NET3 XXOR0.XI1.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI1.XI1.MPMOS1 XXOR0.XI1.NET3 XXOR0.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI2.MNMOS0 XXOR0.XI2.XI2.NET2 XXOR0.XI2.NET2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI2.MNMOS1 NET37 XXOR0.XI2.NET3 XXOR0.XI2.XI2.NET2 VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI2.XI2.MPMOS0 NET37 XXOR0.XI2.NET2 VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07
+ AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI2.MPMOS1 NET37 XXOR0.XI2.NET3 VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07
+ AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI0.MNMOS0 XXOR0.XI2.XI0.NET2 STATE<0> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI0.MNMOS1 XXOR0.XI2.NET2 XXOR0.XI2.NET1 XXOR0.XI2.XI0.NET2 VSS!
+ NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI2.XI0.MPMOS0 XXOR0.XI2.NET2 STATE<0> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI0.MPMOS1 XXOR0.XI2.NET2 XXOR0.XI2.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.Xnand0.MNMOS0 XXOR0.XI2.XNAND0.NET2 STATE<0> VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.Xnand0.MNMOS1 XXOR0.XI2.NET1 XXOR0.NET2 XXOR0.XI2.XNAND0.NET2 VSS!
+ NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI2.Xnand0.MPMOS0 XXOR0.XI2.NET1 STATE<0> VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.Xnand0.MPMOS1 XXOR0.XI2.NET1 XXOR0.NET2 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI1.MNMOS0 XXOR0.XI2.XI1.NET2 XXOR0.XI2.NET1 VSS! VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI1.MNMOS1 XXOR0.XI2.NET3 XXOR0.NET2 XXOR0.XI2.XI1.NET2 VSS! NMOS_VTG
+ L=6e-08 W=3.5e-07 AD=3.675e-14 AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXxor0.XI2.XI1.MPMOS0 XXOR0.XI2.NET3 XXOR0.XI2.NET1 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXxor0.XI2.XI1.MPMOS1 XXOR0.XI2.NET3 XXOR0.NET2 VDD! VDD! PMOS_VTG L=6e-08
+ W=3.5e-07 AD=5.6e-14 AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXor0.XI1.MM0 NET35 XOR0.NET1 VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXor0.XI1.MM1 NET35 XOR0.NET1 VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXor0.XI0.MNMOS0 XOR0.NET1 RST VSS! VSS! NMOS_VTG L=6e-08 W=9.5e-08 AD=1.52e-14
+ AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXor0.XI0.MNMOS1 XOR0.NET1 NET37 VSS! VSS! NMOS_VTG L=6e-08 W=9.5e-08
+ AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXor0.XI0.MPMOS0 XOR0.XI0.NET1 RST VDD! VDD! PMOS_VTG L=6e-08 W=3.55e-07
+ AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXor0.XI0.MPMOS1 XOR0.NET1 NET37 XOR0.XI0.NET1 VDD! PMOS_VTG L=6e-08 W=3.55e-07
+ AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr15.Xml0.Xnand0.MNMOS1 XDFSR15.XML0.XNAND0.NET2 XDFSR15.N VSS! VSS!
+ NMOS_VTG L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr15.Xml0.Xnand0.MNMOS0 XDFSR15.XML0.N4 XDFSR15.RST_BAR
+ XDFSR15.XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14
+ PD=7.1e-07 PS=8.2e-07
mXdfsr15.Xml0.Xnand0.MPMOS1 XDFSR15.XML0.N4 XDFSR15.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr15.Xml0.Xnand0.MPMOS0 XDFSR15.XML0.N4 XDFSR15.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr15.Xml0.Xi0.MM0 XDFSR15.XML0.N1 NET35 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xml0.Xi0.MM1 XDFSR15.XML0.N1 NET35 VDD! VDD! PMOS_VTG L=6e-08 W=4.1e-07
+ AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr15.Xml0.Xi1.MM0 XDFSR15.N XDFSR15.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xml0.Xi1.MM1 XDFSR15.N XDFSR15.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr15.Xsl0.Xi0.MM0 XDFSR15.XSL0.N2 XDFSR15.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xsl0.Xi0.MM1 XDFSR15.XSL0.N2 XDFSR15.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr15.Xsl0.Xi1.MM0 STATE<15> XDFSR15.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xsl0.Xi1.MM1 STATE<15> XDFSR15.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr15.XI0.MM0 XDFSR15.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr15.XI0.MM1 XDFSR15.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr15.XI1.MM0 XDFSR15.CLKI XDFSR15.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr15.XI1.MM1 XDFSR15.CLKI XDFSR15.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr15.XI2.MM0 XDFSR15.RST_BAR VSS! VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr15.XI2.MM1 XDFSR15.RST_BAR VSS! VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr15.Xsl0.Xnor0.MNMOS1 XDFSR15.XSL0.N3 XDFSR15.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr15.Xsl0.Xnor0.MNMOS0 XDFSR15.XSL0.N3 VSS! VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr15.Xsl0.Xnor0.MPMOS1 XDFSR15.XSL0.XNOR0.NET1 XDFSR15.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr15.Xsl0.Xnor0.MPMOS0 XDFSR15.XSL0.N3 VSS! XDFSR15.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr15.Xml0.Xtg0.MM0 XDFSR15.XML0.N1 XDFSR15.CLKI_BAR XDFSR15.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr15.Xml0.Xtg0.MM1 XDFSR15.XML0.N1 XDFSR15.CLKI XDFSR15.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xml0.Xtg1.MM0 XDFSR15.XML0.N4 XDFSR15.CLKI XDFSR15.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr15.Xml0.Xtg1.MM1 XDFSR15.XML0.N4 XDFSR15.CLKI_BAR XDFSR15.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xsl0.Xtg1.MM0 XDFSR15.N XDFSR15.CLKI XDFSR15.XSL0.N1 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr15.Xsl0.Xtg1.MM1 XDFSR15.N XDFSR15.CLKI_BAR XDFSR15.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr15.Xsl0.Xtg0.MM0 XDFSR15.XSL0.N3 XDFSR15.CLKI_BAR XDFSR15.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr15.Xsl0.Xtg0.MM1 XDFSR15.XSL0.N3 XDFSR15.CLKI XDFSR15.XSL0.N1 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xml0.Xnand0.MNMOS1 XDFSR14.XML0.XNAND0.NET2 XDFSR14.N VSS! VSS!
+ NMOS_VTG L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr14.Xml0.Xnand0.MNMOS0 XDFSR14.XML0.N4 XDFSR14.RST_BAR
+ XDFSR14.XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14
+ PD=7.1e-07 PS=8.2e-07
mXdfsr14.Xml0.Xnand0.MPMOS1 XDFSR14.XML0.N4 XDFSR14.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr14.Xml0.Xnand0.MPMOS0 XDFSR14.XML0.N4 XDFSR14.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr14.Xml0.Xi0.MM0 XDFSR14.XML0.N1 STATE<15> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xml0.Xi0.MM1 XDFSR14.XML0.N1 STATE<15> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr14.Xml0.Xi1.MM0 XDFSR14.N XDFSR14.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xml0.Xi1.MM1 XDFSR14.N XDFSR14.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr14.Xsl0.Xi0.MM0 XDFSR14.XSL0.N2 XDFSR14.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xsl0.Xi0.MM1 XDFSR14.XSL0.N2 XDFSR14.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr14.Xsl0.Xi1.MM0 STATE<14> XDFSR14.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xsl0.Xi1.MM1 STATE<14> XDFSR14.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr14.XI0.MM0 XDFSR14.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr14.XI0.MM1 XDFSR14.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr14.XI1.MM0 XDFSR14.CLKI XDFSR14.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr14.XI1.MM1 XDFSR14.CLKI XDFSR14.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr14.XI2.MM0 XDFSR14.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr14.XI2.MM1 XDFSR14.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr14.Xsl0.Xnor0.MNMOS1 XDFSR14.XSL0.N3 XDFSR14.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr14.Xsl0.Xnor0.MNMOS0 XDFSR14.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr14.Xsl0.Xnor0.MPMOS1 XDFSR14.XSL0.XNOR0.NET1 XDFSR14.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr14.Xsl0.Xnor0.MPMOS0 XDFSR14.XSL0.N3 RST XDFSR14.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr14.Xml0.Xtg0.MM0 XDFSR14.XML0.N1 XDFSR14.CLKI_BAR XDFSR14.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr14.Xml0.Xtg0.MM1 XDFSR14.XML0.N1 XDFSR14.CLKI XDFSR14.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xml0.Xtg1.MM0 XDFSR14.XML0.N4 XDFSR14.CLKI XDFSR14.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr14.Xml0.Xtg1.MM1 XDFSR14.XML0.N4 XDFSR14.CLKI_BAR XDFSR14.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xsl0.Xtg1.MM0 XDFSR14.N XDFSR14.CLKI XDFSR14.XSL0.N1 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr14.Xsl0.Xtg1.MM1 XDFSR14.N XDFSR14.CLKI_BAR XDFSR14.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr14.Xsl0.Xtg0.MM0 XDFSR14.XSL0.N3 XDFSR14.CLKI_BAR XDFSR14.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr14.Xsl0.Xtg0.MM1 XDFSR14.XSL0.N3 XDFSR14.CLKI XDFSR14.XSL0.N1 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xml0.Xnand0.MNMOS1 XDFSR13.XML0.XNAND0.NET2 XDFSR13.N VSS! VSS!
+ NMOS_VTG L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr13.Xml0.Xnand0.MNMOS0 XDFSR13.XML0.N4 XDFSR13.RST_BAR
+ XDFSR13.XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14
+ PD=7.1e-07 PS=8.2e-07
mXdfsr13.Xml0.Xnand0.MPMOS1 XDFSR13.XML0.N4 XDFSR13.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr13.Xml0.Xnand0.MPMOS0 XDFSR13.XML0.N4 XDFSR13.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr13.Xml0.Xi0.MM0 XDFSR13.XML0.N1 STATE<14> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xml0.Xi0.MM1 XDFSR13.XML0.N1 STATE<14> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr13.Xml0.Xi1.MM0 XDFSR13.N XDFSR13.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xml0.Xi1.MM1 XDFSR13.N XDFSR13.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr13.Xsl0.Xi0.MM0 XDFSR13.XSL0.N2 XDFSR13.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xsl0.Xi0.MM1 XDFSR13.XSL0.N2 XDFSR13.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr13.Xsl0.Xi1.MM0 STATE<13> XDFSR13.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xsl0.Xi1.MM1 STATE<13> XDFSR13.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr13.XI0.MM0 XDFSR13.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr13.XI0.MM1 XDFSR13.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr13.XI1.MM0 XDFSR13.CLKI XDFSR13.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr13.XI1.MM1 XDFSR13.CLKI XDFSR13.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr13.XI2.MM0 XDFSR13.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr13.XI2.MM1 XDFSR13.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr13.Xsl0.Xnor0.MNMOS1 XDFSR13.XSL0.N3 XDFSR13.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr13.Xsl0.Xnor0.MNMOS0 XDFSR13.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr13.Xsl0.Xnor0.MPMOS1 XDFSR13.XSL0.XNOR0.NET1 XDFSR13.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr13.Xsl0.Xnor0.MPMOS0 XDFSR13.XSL0.N3 RST XDFSR13.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr13.Xml0.Xtg0.MM0 XDFSR13.XML0.N1 XDFSR13.CLKI_BAR XDFSR13.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr13.Xml0.Xtg0.MM1 XDFSR13.XML0.N1 XDFSR13.CLKI XDFSR13.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xml0.Xtg1.MM0 XDFSR13.XML0.N4 XDFSR13.CLKI XDFSR13.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr13.Xml0.Xtg1.MM1 XDFSR13.XML0.N4 XDFSR13.CLKI_BAR XDFSR13.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xsl0.Xtg1.MM0 XDFSR13.N XDFSR13.CLKI XDFSR13.XSL0.N1 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr13.Xsl0.Xtg1.MM1 XDFSR13.N XDFSR13.CLKI_BAR XDFSR13.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr13.Xsl0.Xtg0.MM0 XDFSR13.XSL0.N3 XDFSR13.CLKI_BAR XDFSR13.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr13.Xsl0.Xtg0.MM1 XDFSR13.XSL0.N3 XDFSR13.CLKI XDFSR13.XSL0.N1 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xml0.Xnand0.MNMOS1 XDFSR12.XML0.XNAND0.NET2 XDFSR12.N VSS! VSS!
+ NMOS_VTG L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr12.Xml0.Xnand0.MNMOS0 XDFSR12.XML0.N4 XDFSR12.RST_BAR
+ XDFSR12.XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14
+ PD=7.1e-07 PS=8.2e-07
mXdfsr12.Xml0.Xnand0.MPMOS1 XDFSR12.XML0.N4 XDFSR12.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr12.Xml0.Xnand0.MPMOS0 XDFSR12.XML0.N4 XDFSR12.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr12.Xml0.Xi0.MM0 XDFSR12.XML0.N1 STATE<13> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xml0.Xi0.MM1 XDFSR12.XML0.N1 STATE<13> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr12.Xml0.Xi1.MM0 XDFSR12.N XDFSR12.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xml0.Xi1.MM1 XDFSR12.N XDFSR12.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr12.Xsl0.Xi0.MM0 XDFSR12.XSL0.N2 XDFSR12.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xsl0.Xi0.MM1 XDFSR12.XSL0.N2 XDFSR12.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr12.Xsl0.Xi1.MM0 STATE<12> XDFSR12.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xsl0.Xi1.MM1 STATE<12> XDFSR12.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr12.XI0.MM0 XDFSR12.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr12.XI0.MM1 XDFSR12.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr12.XI1.MM0 XDFSR12.CLKI XDFSR12.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr12.XI1.MM1 XDFSR12.CLKI XDFSR12.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr12.XI2.MM0 XDFSR12.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr12.XI2.MM1 XDFSR12.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr12.Xsl0.Xnor0.MNMOS1 XDFSR12.XSL0.N3 XDFSR12.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr12.Xsl0.Xnor0.MNMOS0 XDFSR12.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr12.Xsl0.Xnor0.MPMOS1 XDFSR12.XSL0.XNOR0.NET1 XDFSR12.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr12.Xsl0.Xnor0.MPMOS0 XDFSR12.XSL0.N3 RST XDFSR12.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr12.Xml0.Xtg0.MM0 XDFSR12.XML0.N1 XDFSR12.CLKI_BAR XDFSR12.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr12.Xml0.Xtg0.MM1 XDFSR12.XML0.N1 XDFSR12.CLKI XDFSR12.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xml0.Xtg1.MM0 XDFSR12.XML0.N4 XDFSR12.CLKI XDFSR12.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr12.Xml0.Xtg1.MM1 XDFSR12.XML0.N4 XDFSR12.CLKI_BAR XDFSR12.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xsl0.Xtg1.MM0 XDFSR12.N XDFSR12.CLKI XDFSR12.XSL0.N1 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr12.Xsl0.Xtg1.MM1 XDFSR12.N XDFSR12.CLKI_BAR XDFSR12.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr12.Xsl0.Xtg0.MM0 XDFSR12.XSL0.N3 XDFSR12.CLKI_BAR XDFSR12.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr12.Xsl0.Xtg0.MM1 XDFSR12.XSL0.N3 XDFSR12.CLKI XDFSR12.XSL0.N1 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xml0.Xnand0.MNMOS1 XDFSR11.XML0.XNAND0.NET2 XDFSR11.N VSS! VSS!
+ NMOS_VTG L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr11.Xml0.Xnand0.MNMOS0 XDFSR11.XML0.N4 XDFSR11.RST_BAR
+ XDFSR11.XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14
+ PD=7.1e-07 PS=8.2e-07
mXdfsr11.Xml0.Xnand0.MPMOS1 XDFSR11.XML0.N4 XDFSR11.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr11.Xml0.Xnand0.MPMOS0 XDFSR11.XML0.N4 XDFSR11.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr11.Xml0.Xi0.MM0 XDFSR11.XML0.N1 STATE<12> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xml0.Xi0.MM1 XDFSR11.XML0.N1 STATE<12> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr11.Xml0.Xi1.MM0 XDFSR11.N XDFSR11.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xml0.Xi1.MM1 XDFSR11.N XDFSR11.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr11.Xsl0.Xi0.MM0 XDFSR11.XSL0.N2 XDFSR11.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xsl0.Xi0.MM1 XDFSR11.XSL0.N2 XDFSR11.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr11.Xsl0.Xi1.MM0 STATE<11> XDFSR11.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xsl0.Xi1.MM1 STATE<11> XDFSR11.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr11.XI0.MM0 XDFSR11.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr11.XI0.MM1 XDFSR11.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr11.XI1.MM0 XDFSR11.CLKI XDFSR11.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr11.XI1.MM1 XDFSR11.CLKI XDFSR11.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr11.XI2.MM0 XDFSR11.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr11.XI2.MM1 XDFSR11.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr11.Xsl0.Xnor0.MNMOS1 XDFSR11.XSL0.N3 XDFSR11.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr11.Xsl0.Xnor0.MNMOS0 XDFSR11.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr11.Xsl0.Xnor0.MPMOS1 XDFSR11.XSL0.XNOR0.NET1 XDFSR11.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr11.Xsl0.Xnor0.MPMOS0 XDFSR11.XSL0.N3 RST XDFSR11.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr11.Xml0.Xtg0.MM0 XDFSR11.XML0.N1 XDFSR11.CLKI_BAR XDFSR11.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr11.Xml0.Xtg0.MM1 XDFSR11.XML0.N1 XDFSR11.CLKI XDFSR11.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xml0.Xtg1.MM0 XDFSR11.XML0.N4 XDFSR11.CLKI XDFSR11.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr11.Xml0.Xtg1.MM1 XDFSR11.XML0.N4 XDFSR11.CLKI_BAR XDFSR11.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xsl0.Xtg1.MM0 XDFSR11.N XDFSR11.CLKI XDFSR11.XSL0.N1 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr11.Xsl0.Xtg1.MM1 XDFSR11.N XDFSR11.CLKI_BAR XDFSR11.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr11.Xsl0.Xtg0.MM0 XDFSR11.XSL0.N3 XDFSR11.CLKI_BAR XDFSR11.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr11.Xsl0.Xtg0.MM1 XDFSR11.XSL0.N3 XDFSR11.CLKI XDFSR11.XSL0.N1 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xml0.Xnand0.MNMOS1 XDFSR10.XML0.XNAND0.NET2 XDFSR10.N VSS! VSS!
+ NMOS_VTG L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr10.Xml0.Xnand0.MNMOS0 XDFSR10.XML0.N4 XDFSR10.RST_BAR
+ XDFSR10.XML0.XNAND0.NET2 VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14
+ PD=7.1e-07 PS=8.2e-07
mXdfsr10.Xml0.Xnand0.MPMOS1 XDFSR10.XML0.N4 XDFSR10.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr10.Xml0.Xnand0.MPMOS0 XDFSR10.XML0.N4 XDFSR10.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr10.Xml0.Xi0.MM0 XDFSR10.XML0.N1 STATE<11> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xml0.Xi0.MM1 XDFSR10.XML0.N1 STATE<11> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr10.Xml0.Xi1.MM0 XDFSR10.N XDFSR10.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xml0.Xi1.MM1 XDFSR10.N XDFSR10.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr10.Xsl0.Xi0.MM0 XDFSR10.XSL0.N2 XDFSR10.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xsl0.Xi0.MM1 XDFSR10.XSL0.N2 XDFSR10.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr10.Xsl0.Xi1.MM0 STATE<10> XDFSR10.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xsl0.Xi1.MM1 STATE<10> XDFSR10.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr10.XI0.MM0 XDFSR10.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr10.XI0.MM1 XDFSR10.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr10.XI1.MM0 XDFSR10.CLKI XDFSR10.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr10.XI1.MM1 XDFSR10.CLKI XDFSR10.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr10.XI2.MM0 XDFSR10.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr10.XI2.MM1 XDFSR10.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr10.Xsl0.Xnor0.MNMOS1 XDFSR10.XSL0.N3 XDFSR10.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr10.Xsl0.Xnor0.MNMOS0 XDFSR10.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr10.Xsl0.Xnor0.MPMOS1 XDFSR10.XSL0.XNOR0.NET1 XDFSR10.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr10.Xsl0.Xnor0.MPMOS0 XDFSR10.XSL0.N3 RST XDFSR10.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr10.Xml0.Xtg0.MM0 XDFSR10.XML0.N1 XDFSR10.CLKI_BAR XDFSR10.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr10.Xml0.Xtg0.MM1 XDFSR10.XML0.N1 XDFSR10.CLKI XDFSR10.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xml0.Xtg1.MM0 XDFSR10.XML0.N4 XDFSR10.CLKI XDFSR10.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr10.Xml0.Xtg1.MM1 XDFSR10.XML0.N4 XDFSR10.CLKI_BAR XDFSR10.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xsl0.Xtg1.MM0 XDFSR10.N XDFSR10.CLKI XDFSR10.XSL0.N1 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr10.Xsl0.Xtg1.MM1 XDFSR10.N XDFSR10.CLKI_BAR XDFSR10.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr10.Xsl0.Xtg0.MM0 XDFSR10.XSL0.N3 XDFSR10.CLKI_BAR XDFSR10.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr10.Xsl0.Xtg0.MM1 XDFSR10.XSL0.N3 XDFSR10.CLKI XDFSR10.XSL0.N1 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xml0.Xnand0.MNMOS1 XDFSR9.XML0.XNAND0.NET2 XDFSR9.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr9.Xml0.Xnand0.MNMOS0 XDFSR9.XML0.N4 XDFSR9.RST_BAR XDFSR9.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr9.Xml0.Xnand0.MPMOS1 XDFSR9.XML0.N4 XDFSR9.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr9.Xml0.Xnand0.MPMOS0 XDFSR9.XML0.N4 XDFSR9.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr9.Xml0.Xi0.MM0 XDFSR9.XML0.N1 STATE<10> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xml0.Xi0.MM1 XDFSR9.XML0.N1 STATE<10> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr9.Xml0.Xi1.MM0 XDFSR9.N XDFSR9.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xml0.Xi1.MM1 XDFSR9.N XDFSR9.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr9.Xsl0.Xi0.MM0 XDFSR9.XSL0.N2 XDFSR9.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xsl0.Xi0.MM1 XDFSR9.XSL0.N2 XDFSR9.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr9.Xsl0.Xi1.MM0 STATE<9> XDFSR9.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xsl0.Xi1.MM1 STATE<9> XDFSR9.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr9.XI0.MM0 XDFSR9.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr9.XI0.MM1 XDFSR9.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr9.XI1.MM0 XDFSR9.CLKI XDFSR9.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr9.XI1.MM1 XDFSR9.CLKI XDFSR9.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr9.XI2.MM0 XDFSR9.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr9.XI2.MM1 XDFSR9.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr9.Xsl0.Xnor0.MNMOS1 XDFSR9.XSL0.N3 XDFSR9.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr9.Xsl0.Xnor0.MNMOS0 XDFSR9.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr9.Xsl0.Xnor0.MPMOS1 XDFSR9.XSL0.XNOR0.NET1 XDFSR9.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr9.Xsl0.Xnor0.MPMOS0 XDFSR9.XSL0.N3 RST XDFSR9.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr9.Xml0.Xtg0.MM0 XDFSR9.XML0.N1 XDFSR9.CLKI_BAR XDFSR9.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr9.Xml0.Xtg0.MM1 XDFSR9.XML0.N1 XDFSR9.CLKI XDFSR9.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xml0.Xtg1.MM0 XDFSR9.XML0.N4 XDFSR9.CLKI XDFSR9.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr9.Xml0.Xtg1.MM1 XDFSR9.XML0.N4 XDFSR9.CLKI_BAR XDFSR9.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xsl0.Xtg1.MM0 XDFSR9.N XDFSR9.CLKI XDFSR9.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr9.Xsl0.Xtg1.MM1 XDFSR9.N XDFSR9.CLKI_BAR XDFSR9.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr9.Xsl0.Xtg0.MM0 XDFSR9.XSL0.N3 XDFSR9.CLKI_BAR XDFSR9.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr9.Xsl0.Xtg0.MM1 XDFSR9.XSL0.N3 XDFSR9.CLKI XDFSR9.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xml0.Xnand0.MNMOS1 XDFSR8.XML0.XNAND0.NET2 XDFSR8.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr8.Xml0.Xnand0.MNMOS0 XDFSR8.XML0.N4 XDFSR8.RST_BAR XDFSR8.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr8.Xml0.Xnand0.MPMOS1 XDFSR8.XML0.N4 XDFSR8.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr8.Xml0.Xnand0.MPMOS0 XDFSR8.XML0.N4 XDFSR8.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr8.Xml0.Xi0.MM0 XDFSR8.XML0.N1 STATE<9> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xml0.Xi0.MM1 XDFSR8.XML0.N1 STATE<9> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr8.Xml0.Xi1.MM0 XDFSR8.N XDFSR8.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xml0.Xi1.MM1 XDFSR8.N XDFSR8.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr8.Xsl0.Xi0.MM0 XDFSR8.XSL0.N2 XDFSR8.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xsl0.Xi0.MM1 XDFSR8.XSL0.N2 XDFSR8.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr8.Xsl0.Xi1.MM0 STATE<8> XDFSR8.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xsl0.Xi1.MM1 STATE<8> XDFSR8.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr8.XI0.MM0 XDFSR8.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr8.XI0.MM1 XDFSR8.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr8.XI1.MM0 XDFSR8.CLKI XDFSR8.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr8.XI1.MM1 XDFSR8.CLKI XDFSR8.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr8.XI2.MM0 XDFSR8.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr8.XI2.MM1 XDFSR8.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr8.Xsl0.Xnor0.MNMOS1 XDFSR8.XSL0.N3 XDFSR8.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr8.Xsl0.Xnor0.MNMOS0 XDFSR8.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr8.Xsl0.Xnor0.MPMOS1 XDFSR8.XSL0.XNOR0.NET1 XDFSR8.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr8.Xsl0.Xnor0.MPMOS0 XDFSR8.XSL0.N3 RST XDFSR8.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr8.Xml0.Xtg0.MM0 XDFSR8.XML0.N1 XDFSR8.CLKI_BAR XDFSR8.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr8.Xml0.Xtg0.MM1 XDFSR8.XML0.N1 XDFSR8.CLKI XDFSR8.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xml0.Xtg1.MM0 XDFSR8.XML0.N4 XDFSR8.CLKI XDFSR8.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr8.Xml0.Xtg1.MM1 XDFSR8.XML0.N4 XDFSR8.CLKI_BAR XDFSR8.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xsl0.Xtg1.MM0 XDFSR8.N XDFSR8.CLKI XDFSR8.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr8.Xsl0.Xtg1.MM1 XDFSR8.N XDFSR8.CLKI_BAR XDFSR8.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr8.Xsl0.Xtg0.MM0 XDFSR8.XSL0.N3 XDFSR8.CLKI_BAR XDFSR8.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr8.Xsl0.Xtg0.MM1 XDFSR8.XSL0.N3 XDFSR8.CLKI XDFSR8.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xml0.Xnand0.MNMOS1 XDFSR7.XML0.XNAND0.NET2 XDFSR7.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr7.Xml0.Xnand0.MNMOS0 XDFSR7.XML0.N4 XDFSR7.RST_BAR XDFSR7.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr7.Xml0.Xnand0.MPMOS1 XDFSR7.XML0.N4 XDFSR7.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr7.Xml0.Xnand0.MPMOS0 XDFSR7.XML0.N4 XDFSR7.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr7.Xml0.Xi0.MM0 XDFSR7.XML0.N1 STATE<8> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xml0.Xi0.MM1 XDFSR7.XML0.N1 STATE<8> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr7.Xml0.Xi1.MM0 XDFSR7.N XDFSR7.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xml0.Xi1.MM1 XDFSR7.N XDFSR7.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr7.Xsl0.Xi0.MM0 XDFSR7.XSL0.N2 XDFSR7.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xsl0.Xi0.MM1 XDFSR7.XSL0.N2 XDFSR7.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr7.Xsl0.Xi1.MM0 STATE<7> XDFSR7.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xsl0.Xi1.MM1 STATE<7> XDFSR7.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr7.XI0.MM0 XDFSR7.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr7.XI0.MM1 XDFSR7.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr7.XI1.MM0 XDFSR7.CLKI XDFSR7.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr7.XI1.MM1 XDFSR7.CLKI XDFSR7.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr7.XI2.MM0 XDFSR7.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr7.XI2.MM1 XDFSR7.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr7.Xsl0.Xnor0.MNMOS1 XDFSR7.XSL0.N3 XDFSR7.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr7.Xsl0.Xnor0.MNMOS0 XDFSR7.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr7.Xsl0.Xnor0.MPMOS1 XDFSR7.XSL0.XNOR0.NET1 XDFSR7.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr7.Xsl0.Xnor0.MPMOS0 XDFSR7.XSL0.N3 RST XDFSR7.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr7.Xml0.Xtg0.MM0 XDFSR7.XML0.N1 XDFSR7.CLKI_BAR XDFSR7.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr7.Xml0.Xtg0.MM1 XDFSR7.XML0.N1 XDFSR7.CLKI XDFSR7.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xml0.Xtg1.MM0 XDFSR7.XML0.N4 XDFSR7.CLKI XDFSR7.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr7.Xml0.Xtg1.MM1 XDFSR7.XML0.N4 XDFSR7.CLKI_BAR XDFSR7.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xsl0.Xtg1.MM0 XDFSR7.N XDFSR7.CLKI XDFSR7.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr7.Xsl0.Xtg1.MM1 XDFSR7.N XDFSR7.CLKI_BAR XDFSR7.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr7.Xsl0.Xtg0.MM0 XDFSR7.XSL0.N3 XDFSR7.CLKI_BAR XDFSR7.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr7.Xsl0.Xtg0.MM1 XDFSR7.XSL0.N3 XDFSR7.CLKI XDFSR7.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xml0.Xnand0.MNMOS1 XDFSR6.XML0.XNAND0.NET2 XDFSR6.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr6.Xml0.Xnand0.MNMOS0 XDFSR6.XML0.N4 XDFSR6.RST_BAR XDFSR6.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr6.Xml0.Xnand0.MPMOS1 XDFSR6.XML0.N4 XDFSR6.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr6.Xml0.Xnand0.MPMOS0 XDFSR6.XML0.N4 XDFSR6.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr6.Xml0.Xi0.MM0 XDFSR6.XML0.N1 STATE<7> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xml0.Xi0.MM1 XDFSR6.XML0.N1 STATE<7> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr6.Xml0.Xi1.MM0 XDFSR6.N XDFSR6.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xml0.Xi1.MM1 XDFSR6.N XDFSR6.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr6.Xsl0.Xi0.MM0 XDFSR6.XSL0.N2 XDFSR6.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xsl0.Xi0.MM1 XDFSR6.XSL0.N2 XDFSR6.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr6.Xsl0.Xi1.MM0 STATE<6> XDFSR6.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xsl0.Xi1.MM1 STATE<6> XDFSR6.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr6.XI0.MM0 XDFSR6.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr6.XI0.MM1 XDFSR6.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr6.XI1.MM0 XDFSR6.CLKI XDFSR6.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr6.XI1.MM1 XDFSR6.CLKI XDFSR6.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr6.XI2.MM0 XDFSR6.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr6.XI2.MM1 XDFSR6.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr6.Xsl0.Xnor0.MNMOS1 XDFSR6.XSL0.N3 XDFSR6.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr6.Xsl0.Xnor0.MNMOS0 XDFSR6.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr6.Xsl0.Xnor0.MPMOS1 XDFSR6.XSL0.XNOR0.NET1 XDFSR6.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr6.Xsl0.Xnor0.MPMOS0 XDFSR6.XSL0.N3 RST XDFSR6.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr6.Xml0.Xtg0.MM0 XDFSR6.XML0.N1 XDFSR6.CLKI_BAR XDFSR6.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr6.Xml0.Xtg0.MM1 XDFSR6.XML0.N1 XDFSR6.CLKI XDFSR6.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xml0.Xtg1.MM0 XDFSR6.XML0.N4 XDFSR6.CLKI XDFSR6.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr6.Xml0.Xtg1.MM1 XDFSR6.XML0.N4 XDFSR6.CLKI_BAR XDFSR6.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xsl0.Xtg1.MM0 XDFSR6.N XDFSR6.CLKI XDFSR6.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr6.Xsl0.Xtg1.MM1 XDFSR6.N XDFSR6.CLKI_BAR XDFSR6.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr6.Xsl0.Xtg0.MM0 XDFSR6.XSL0.N3 XDFSR6.CLKI_BAR XDFSR6.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr6.Xsl0.Xtg0.MM1 XDFSR6.XSL0.N3 XDFSR6.CLKI XDFSR6.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xml0.Xnand0.MNMOS1 XDFSR5.XML0.XNAND0.NET2 XDFSR5.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr5.Xml0.Xnand0.MNMOS0 XDFSR5.XML0.N4 XDFSR5.RST_BAR XDFSR5.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr5.Xml0.Xnand0.MPMOS1 XDFSR5.XML0.N4 XDFSR5.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr5.Xml0.Xnand0.MPMOS0 XDFSR5.XML0.N4 XDFSR5.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr5.Xml0.Xi0.MM0 XDFSR5.XML0.N1 STATE<6> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xml0.Xi0.MM1 XDFSR5.XML0.N1 STATE<6> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr5.Xml0.Xi1.MM0 XDFSR5.N XDFSR5.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xml0.Xi1.MM1 XDFSR5.N XDFSR5.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr5.Xsl0.Xi0.MM0 XDFSR5.XSL0.N2 XDFSR5.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xsl0.Xi0.MM1 XDFSR5.XSL0.N2 XDFSR5.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr5.Xsl0.Xi1.MM0 STATE<5> XDFSR5.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xsl0.Xi1.MM1 STATE<5> XDFSR5.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr5.XI0.MM0 XDFSR5.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr5.XI0.MM1 XDFSR5.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr5.XI1.MM0 XDFSR5.CLKI XDFSR5.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr5.XI1.MM1 XDFSR5.CLKI XDFSR5.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr5.XI2.MM0 XDFSR5.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr5.XI2.MM1 XDFSR5.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr5.Xsl0.Xnor0.MNMOS1 XDFSR5.XSL0.N3 XDFSR5.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr5.Xsl0.Xnor0.MNMOS0 XDFSR5.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr5.Xsl0.Xnor0.MPMOS1 XDFSR5.XSL0.XNOR0.NET1 XDFSR5.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr5.Xsl0.Xnor0.MPMOS0 XDFSR5.XSL0.N3 RST XDFSR5.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr5.Xml0.Xtg0.MM0 XDFSR5.XML0.N1 XDFSR5.CLKI_BAR XDFSR5.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr5.Xml0.Xtg0.MM1 XDFSR5.XML0.N1 XDFSR5.CLKI XDFSR5.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xml0.Xtg1.MM0 XDFSR5.XML0.N4 XDFSR5.CLKI XDFSR5.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr5.Xml0.Xtg1.MM1 XDFSR5.XML0.N4 XDFSR5.CLKI_BAR XDFSR5.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xsl0.Xtg1.MM0 XDFSR5.N XDFSR5.CLKI XDFSR5.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr5.Xsl0.Xtg1.MM1 XDFSR5.N XDFSR5.CLKI_BAR XDFSR5.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr5.Xsl0.Xtg0.MM0 XDFSR5.XSL0.N3 XDFSR5.CLKI_BAR XDFSR5.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr5.Xsl0.Xtg0.MM1 XDFSR5.XSL0.N3 XDFSR5.CLKI XDFSR5.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xml0.Xnand0.MNMOS1 XDFSR4.XML0.XNAND0.NET2 XDFSR4.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr4.Xml0.Xnand0.MNMOS0 XDFSR4.XML0.N4 XDFSR4.RST_BAR XDFSR4.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr4.Xml0.Xnand0.MPMOS1 XDFSR4.XML0.N4 XDFSR4.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr4.Xml0.Xnand0.MPMOS0 XDFSR4.XML0.N4 XDFSR4.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr4.Xml0.Xi0.MM0 XDFSR4.XML0.N1 STATE<5> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xml0.Xi0.MM1 XDFSR4.XML0.N1 STATE<5> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr4.Xml0.Xi1.MM0 XDFSR4.N XDFSR4.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xml0.Xi1.MM1 XDFSR4.N XDFSR4.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr4.Xsl0.Xi0.MM0 XDFSR4.XSL0.N2 XDFSR4.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xsl0.Xi0.MM1 XDFSR4.XSL0.N2 XDFSR4.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr4.Xsl0.Xi1.MM0 STATE<4> XDFSR4.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xsl0.Xi1.MM1 STATE<4> XDFSR4.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr4.XI0.MM0 XDFSR4.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr4.XI0.MM1 XDFSR4.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr4.XI1.MM0 XDFSR4.CLKI XDFSR4.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr4.XI1.MM1 XDFSR4.CLKI XDFSR4.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr4.XI2.MM0 XDFSR4.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr4.XI2.MM1 XDFSR4.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr4.Xsl0.Xnor0.MNMOS1 XDFSR4.XSL0.N3 XDFSR4.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr4.Xsl0.Xnor0.MNMOS0 XDFSR4.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr4.Xsl0.Xnor0.MPMOS1 XDFSR4.XSL0.XNOR0.NET1 XDFSR4.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr4.Xsl0.Xnor0.MPMOS0 XDFSR4.XSL0.N3 RST XDFSR4.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr4.Xml0.Xtg0.MM0 XDFSR4.XML0.N1 XDFSR4.CLKI_BAR XDFSR4.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr4.Xml0.Xtg0.MM1 XDFSR4.XML0.N1 XDFSR4.CLKI XDFSR4.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xml0.Xtg1.MM0 XDFSR4.XML0.N4 XDFSR4.CLKI XDFSR4.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr4.Xml0.Xtg1.MM1 XDFSR4.XML0.N4 XDFSR4.CLKI_BAR XDFSR4.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xsl0.Xtg1.MM0 XDFSR4.N XDFSR4.CLKI XDFSR4.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr4.Xsl0.Xtg1.MM1 XDFSR4.N XDFSR4.CLKI_BAR XDFSR4.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr4.Xsl0.Xtg0.MM0 XDFSR4.XSL0.N3 XDFSR4.CLKI_BAR XDFSR4.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr4.Xsl0.Xtg0.MM1 XDFSR4.XSL0.N3 XDFSR4.CLKI XDFSR4.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xml0.Xnand0.MNMOS1 XDFSR3.XML0.XNAND0.NET2 XDFSR3.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr3.Xml0.Xnand0.MNMOS0 XDFSR3.XML0.N4 XDFSR3.RST_BAR XDFSR3.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr3.Xml0.Xnand0.MPMOS1 XDFSR3.XML0.N4 XDFSR3.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr3.Xml0.Xnand0.MPMOS0 XDFSR3.XML0.N4 XDFSR3.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr3.Xml0.Xi0.MM0 XDFSR3.XML0.N1 STATE<4> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xml0.Xi0.MM1 XDFSR3.XML0.N1 STATE<4> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr3.Xml0.Xi1.MM0 XDFSR3.N XDFSR3.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xml0.Xi1.MM1 XDFSR3.N XDFSR3.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr3.Xsl0.Xi0.MM0 XDFSR3.XSL0.N2 XDFSR3.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xsl0.Xi0.MM1 XDFSR3.XSL0.N2 XDFSR3.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr3.Xsl0.Xi1.MM0 STATE<3> XDFSR3.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xsl0.Xi1.MM1 STATE<3> XDFSR3.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr3.XI0.MM0 XDFSR3.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr3.XI0.MM1 XDFSR3.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr3.XI1.MM0 XDFSR3.CLKI XDFSR3.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr3.XI1.MM1 XDFSR3.CLKI XDFSR3.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr3.XI2.MM0 XDFSR3.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr3.XI2.MM1 XDFSR3.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr3.Xsl0.Xnor0.MNMOS1 XDFSR3.XSL0.N3 XDFSR3.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr3.Xsl0.Xnor0.MNMOS0 XDFSR3.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr3.Xsl0.Xnor0.MPMOS1 XDFSR3.XSL0.XNOR0.NET1 XDFSR3.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr3.Xsl0.Xnor0.MPMOS0 XDFSR3.XSL0.N3 RST XDFSR3.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr3.Xml0.Xtg0.MM0 XDFSR3.XML0.N1 XDFSR3.CLKI_BAR XDFSR3.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr3.Xml0.Xtg0.MM1 XDFSR3.XML0.N1 XDFSR3.CLKI XDFSR3.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xml0.Xtg1.MM0 XDFSR3.XML0.N4 XDFSR3.CLKI XDFSR3.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr3.Xml0.Xtg1.MM1 XDFSR3.XML0.N4 XDFSR3.CLKI_BAR XDFSR3.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xsl0.Xtg1.MM0 XDFSR3.N XDFSR3.CLKI XDFSR3.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr3.Xsl0.Xtg1.MM1 XDFSR3.N XDFSR3.CLKI_BAR XDFSR3.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr3.Xsl0.Xtg0.MM0 XDFSR3.XSL0.N3 XDFSR3.CLKI_BAR XDFSR3.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr3.Xsl0.Xtg0.MM1 XDFSR3.XSL0.N3 XDFSR3.CLKI XDFSR3.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xml0.Xnand0.MNMOS1 XDFSR2.XML0.XNAND0.NET2 XDFSR2.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr2.Xml0.Xnand0.MNMOS0 XDFSR2.XML0.N4 XDFSR2.RST_BAR XDFSR2.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr2.Xml0.Xnand0.MPMOS1 XDFSR2.XML0.N4 XDFSR2.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr2.Xml0.Xnand0.MPMOS0 XDFSR2.XML0.N4 XDFSR2.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr2.Xml0.Xi0.MM0 XDFSR2.XML0.N1 STATE<3> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xml0.Xi0.MM1 XDFSR2.XML0.N1 STATE<3> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr2.Xml0.Xi1.MM0 XDFSR2.N XDFSR2.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xml0.Xi1.MM1 XDFSR2.N XDFSR2.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr2.Xsl0.Xi0.MM0 XDFSR2.XSL0.N2 XDFSR2.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xsl0.Xi0.MM1 XDFSR2.XSL0.N2 XDFSR2.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr2.Xsl0.Xi1.MM0 STATE<2> XDFSR2.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xsl0.Xi1.MM1 STATE<2> XDFSR2.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr2.XI0.MM0 XDFSR2.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr2.XI0.MM1 XDFSR2.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr2.XI1.MM0 XDFSR2.CLKI XDFSR2.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr2.XI1.MM1 XDFSR2.CLKI XDFSR2.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr2.XI2.MM0 XDFSR2.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr2.XI2.MM1 XDFSR2.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr2.Xsl0.Xnor0.MNMOS1 XDFSR2.XSL0.N3 XDFSR2.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr2.Xsl0.Xnor0.MNMOS0 XDFSR2.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr2.Xsl0.Xnor0.MPMOS1 XDFSR2.XSL0.XNOR0.NET1 XDFSR2.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr2.Xsl0.Xnor0.MPMOS0 XDFSR2.XSL0.N3 RST XDFSR2.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr2.Xml0.Xtg0.MM0 XDFSR2.XML0.N1 XDFSR2.CLKI_BAR XDFSR2.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr2.Xml0.Xtg0.MM1 XDFSR2.XML0.N1 XDFSR2.CLKI XDFSR2.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xml0.Xtg1.MM0 XDFSR2.XML0.N4 XDFSR2.CLKI XDFSR2.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr2.Xml0.Xtg1.MM1 XDFSR2.XML0.N4 XDFSR2.CLKI_BAR XDFSR2.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xsl0.Xtg1.MM0 XDFSR2.N XDFSR2.CLKI XDFSR2.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr2.Xsl0.Xtg1.MM1 XDFSR2.N XDFSR2.CLKI_BAR XDFSR2.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr2.Xsl0.Xtg0.MM0 XDFSR2.XSL0.N3 XDFSR2.CLKI_BAR XDFSR2.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr2.Xsl0.Xtg0.MM1 XDFSR2.XSL0.N3 XDFSR2.CLKI XDFSR2.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xml0.Xnand0.MNMOS1 XDFSR1.XML0.XNAND0.NET2 XDFSR1.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr1.Xml0.Xnand0.MNMOS0 XDFSR1.XML0.N4 XDFSR1.RST_BAR XDFSR1.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr1.Xml0.Xnand0.MPMOS1 XDFSR1.XML0.N4 XDFSR1.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr1.Xml0.Xnand0.MPMOS0 XDFSR1.XML0.N4 XDFSR1.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr1.Xml0.Xi0.MM0 XDFSR1.XML0.N1 STATE<2> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xml0.Xi0.MM1 XDFSR1.XML0.N1 STATE<2> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr1.Xml0.Xi1.MM0 XDFSR1.N XDFSR1.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xml0.Xi1.MM1 XDFSR1.N XDFSR1.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr1.Xsl0.Xi0.MM0 XDFSR1.XSL0.N2 XDFSR1.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xsl0.Xi0.MM1 XDFSR1.XSL0.N2 XDFSR1.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr1.Xsl0.Xi1.MM0 STATE<1> XDFSR1.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xsl0.Xi1.MM1 STATE<1> XDFSR1.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr1.XI0.MM0 XDFSR1.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr1.XI0.MM1 XDFSR1.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr1.XI1.MM0 XDFSR1.CLKI XDFSR1.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr1.XI1.MM1 XDFSR1.CLKI XDFSR1.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr1.XI2.MM0 XDFSR1.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr1.XI2.MM1 XDFSR1.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr1.Xsl0.Xnor0.MNMOS1 XDFSR1.XSL0.N3 XDFSR1.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr1.Xsl0.Xnor0.MNMOS0 XDFSR1.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr1.Xsl0.Xnor0.MPMOS1 XDFSR1.XSL0.XNOR0.NET1 XDFSR1.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr1.Xsl0.Xnor0.MPMOS0 XDFSR1.XSL0.N3 RST XDFSR1.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr1.Xml0.Xtg0.MM0 XDFSR1.XML0.N1 XDFSR1.CLKI_BAR XDFSR1.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr1.Xml0.Xtg0.MM1 XDFSR1.XML0.N1 XDFSR1.CLKI XDFSR1.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xml0.Xtg1.MM0 XDFSR1.XML0.N4 XDFSR1.CLKI XDFSR1.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr1.Xml0.Xtg1.MM1 XDFSR1.XML0.N4 XDFSR1.CLKI_BAR XDFSR1.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xsl0.Xtg1.MM0 XDFSR1.N XDFSR1.CLKI XDFSR1.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr1.Xsl0.Xtg1.MM1 XDFSR1.N XDFSR1.CLKI_BAR XDFSR1.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr1.Xsl0.Xtg0.MM0 XDFSR1.XSL0.N3 XDFSR1.CLKI_BAR XDFSR1.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr1.Xsl0.Xtg0.MM1 XDFSR1.XSL0.N3 XDFSR1.CLKI XDFSR1.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xml0.Xnand0.MNMOS1 XDFSR0.XML0.XNAND0.NET2 XDFSR0.N VSS! VSS! NMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4e-14 AS=2.625e-14 PD=8.2e-07 PS=7.1e-07
mXdfsr0.Xml0.Xnand0.MNMOS0 XDFSR0.XML0.N4 XDFSR0.RST_BAR XDFSR0.XML0.XNAND0.NET2
+ VSS! NMOS_VTG L=6e-08 W=2.5e-07 AD=2.625e-14 AS=4e-14 PD=7.1e-07 PS=8.2e-07
mXdfsr0.Xml0.Xnand0.MPMOS1 XDFSR0.XML0.N4 XDFSR0.N VDD! VDD! PMOS_VTG L=6e-08
+ W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr0.Xml0.Xnand0.MPMOS0 XDFSR0.XML0.N4 XDFSR0.RST_BAR VDD! VDD! PMOS_VTG
+ L=6e-08 W=5.25e-07 AD=8.4e-14 AS=5.5125e-14 PD=1.37e-06 PS=1.26e-06
mXdfsr0.Xml0.Xi0.MM0 XDFSR0.XML0.N1 STATE<1> VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xml0.Xi0.MM1 XDFSR0.XML0.N1 STATE<1> VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr0.Xml0.Xi1.MM0 XDFSR0.N XDFSR0.XML0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xml0.Xi1.MM1 XDFSR0.N XDFSR0.XML0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr0.Xsl0.Xi0.MM0 XDFSR0.XSL0.N2 XDFSR0.XSL0.N1 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xsl0.Xi0.MM1 XDFSR0.XSL0.N2 XDFSR0.XSL0.N1 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr0.Xsl0.Xi1.MM0 STATE<0> XDFSR0.XSL0.N2 VSS! VSS! NMOS_VTG L=6e-08
+ W=3.25e-07 AD=3.4125e-14 AS=3.4125e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xsl0.Xi1.MM1 STATE<0> XDFSR0.XSL0.N2 VDD! VDD! PMOS_VTG L=6e-08
+ W=4.1e-07 AD=4.305e-14 AS=4.305e-14 PD=1.03e-06 PS=1.03e-06
mXdfsr0.XI0.MM0 XDFSR0.CLKI_BAR CLK VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr0.XI0.MM1 XDFSR0.CLKI_BAR CLK VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr0.XI1.MM0 XDFSR0.CLKI XDFSR0.CLKI_BAR VSS! VSS! NMOS_VTG L=6e-08
+ W=3.45e-07 AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr0.XI1.MM1 XDFSR0.CLKI XDFSR0.CLKI_BAR VDD! VDD! PMOS_VTG L=6e-08
+ W=4.35e-07 AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr0.XI2.MM0 XDFSR0.RST_BAR RST VSS! VSS! NMOS_VTG L=6e-08 W=3.45e-07
+ AD=3.6225e-14 AS=3.6225e-14 PD=9e-07 PS=9e-07
mXdfsr0.XI2.MM1 XDFSR0.RST_BAR RST VDD! VDD! PMOS_VTG L=6e-08 W=4.35e-07
+ AD=4.5675e-14 AS=4.5675e-14 PD=1.08e-06 PS=1.08e-06
mXdfsr0.Xsl0.Xnor0.MNMOS1 XDFSR0.XSL0.N3 XDFSR0.XSL0.N2 VSS! VSS! NMOS_VTG
+ L=6e-08 W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr0.Xsl0.Xnor0.MNMOS0 XDFSR0.XSL0.N3 RST VSS! VSS! NMOS_VTG L=6e-08
+ W=9.5e-08 AD=1.52e-14 AS=9.975e-15 PD=5.1e-07 PS=4e-07
mXdfsr0.Xsl0.Xnor0.MPMOS1 XDFSR0.XSL0.XNOR0.NET1 XDFSR0.XSL0.N2 VDD! VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=5.68e-14 AS=3.7275e-14 PD=1.03e-06 PS=9.2e-07
mXdfsr0.Xsl0.Xnor0.MPMOS0 XDFSR0.XSL0.N3 RST XDFSR0.XSL0.XNOR0.NET1 VDD!
+ PMOS_VTG L=6e-08 W=3.55e-07 AD=3.7275e-14 AS=5.68e-14 PD=9.2e-07 PS=1.03e-06
mXdfsr0.Xml0.Xtg0.MM0 XDFSR0.XML0.N1 XDFSR0.CLKI_BAR XDFSR0.XML0.N2 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr0.Xml0.Xtg0.MM1 XDFSR0.XML0.N1 XDFSR0.CLKI XDFSR0.XML0.N2 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xml0.Xtg1.MM0 XDFSR0.XML0.N4 XDFSR0.CLKI XDFSR0.XML0.N2 VSS! NMOS_VTG
+ L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr0.Xml0.Xtg1.MM1 XDFSR0.XML0.N4 XDFSR0.CLKI_BAR XDFSR0.XML0.N2 VDD!
+ PMOS_VTG L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xsl0.Xtg1.MM0 XDFSR0.N XDFSR0.CLKI XDFSR0.XSL0.N1 VSS! NMOS_VTG L=6e-08
+ W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr0.Xsl0.Xtg1.MM1 XDFSR0.N XDFSR0.CLKI_BAR XDFSR0.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
mXdfsr0.Xsl0.Xtg0.MM0 XDFSR0.XSL0.N3 XDFSR0.CLKI_BAR XDFSR0.XSL0.N1 VSS!
+ NMOS_VTG L=6e-08 W=2.65e-07 AD=4.77e-14 AS=4.77e-14 PD=8.9e-07 PS=8.9e-07
mXdfsr0.Xsl0.Xtg0.MM1 XDFSR0.XSL0.N3 XDFSR0.CLKI XDFSR0.XSL0.N1 VDD! PMOS_VTG
+ L=6e-08 W=2.5e-07 AD=4.5e-14 AS=4.5e-14 PD=8.6e-07 PS=8.6e-07
c_98 RST 0 4.86758f
c_292 VSS! 0 5.27622f
c_357 STATE<5> 0 0.983993f
c_396 STATE<2> 0 0.498093f
c_590 VDD! 0 11.8914f
c_599 XOR0.NET1 0 0.12011f
c_609 STATE<15> 0 0.133475f
c_620 STATE<14> 0 0.133475f
c_631 STATE<13> 0 0.133475f
c_642 STATE<12> 0 0.133475f
c_653 STATE<11> 0 0.133475f
c_664 STATE<10> 0 0.133475f
c_675 STATE<9> 0 0.133475f
c_686 STATE<8> 0 0.133475f
c_697 STATE<7> 0 0.133475f
c_708 STATE<6> 0 0.133475f
c_720 STATE<4> 0 0.132127f
c_765 STATE<3> 0 0.462979f
c_779 STATE<1> 0 0.129638f
c_835 NET37 0 2.4659f
c_846 NET35 0 0.161767f
c_865 STATE<0> 0 0.422018f
c_874 XXOR0.NET1 0 0.187825f
c_883 XXOR0.NET2 0 0.191081f
c_952 CLK 0 3.49622f
c_964 XXOR0.XI0.NET3 0 0.145563f
c_976 XXOR0.XI0.NET1 0 0.188265f
c_985 XXOR0.XI0.NET2 0 0.0968779f
c_996 XXOR0.XI1.NET3 0 0.157887f
c_1006 XXOR0.XI1.NET1 0 0.20099f
c_1014 XXOR0.XI1.NET2 0 0.101231f
c_1023 XXOR0.XI2.NET3 0 0.153209f
c_1032 XXOR0.XI2.NET1 0 0.198558f
c_1039 XXOR0.XI2.NET2 0 0.096359f
c_1049 XDFSR15.N 0 0.157125f
c_1064 XDFSR15.RST_BAR 0 0.187903f
c_1079 XDFSR15.CLKI_BAR 0 0.34845f
c_1086 XDFSR15.XML0.N1 0 0.0358798f
c_1095 XDFSR15.XML0.N2 0 0.120116f
c_1104 XDFSR15.XML0.N4 0 0.0454161f
c_1113 XDFSR15.XSL0.N1 0 0.122357f
c_1129 XDFSR15.CLKI 0 0.289564f
c_1138 XDFSR15.XSL0.N2 0 0.190162f
c_1147 XDFSR15.XSL0.N3 0 0.0472116f
c_1156 XDFSR14.N 0 0.157317f
c_1171 XDFSR14.RST_BAR 0 0.187903f
c_1188 XDFSR14.CLKI_BAR 0 0.35929f
c_1195 XDFSR14.XML0.N1 0 0.0363245f
c_1203 XDFSR14.XML0.N2 0 0.123269f
c_1211 XDFSR14.XML0.N4 0 0.0453169f
c_1220 XDFSR14.XSL0.N1 0 0.12236f
c_1236 XDFSR14.CLKI 0 0.30462f
c_1246 XDFSR14.XSL0.N2 0 0.190162f
c_1256 XDFSR14.XSL0.N3 0 0.0472116f
c_1265 XDFSR13.N 0 0.157317f
c_1280 XDFSR13.RST_BAR 0 0.187903f
c_1297 XDFSR13.CLKI_BAR 0 0.35929f
c_1304 XDFSR13.XML0.N1 0 0.0363245f
c_1312 XDFSR13.XML0.N2 0 0.123269f
c_1320 XDFSR13.XML0.N4 0 0.0453169f
c_1329 XDFSR13.XSL0.N1 0 0.12236f
c_1345 XDFSR13.CLKI 0 0.30462f
c_1355 XDFSR13.XSL0.N2 0 0.190162f
c_1365 XDFSR13.XSL0.N3 0 0.0472116f
c_1374 XDFSR12.N 0 0.157317f
c_1389 XDFSR12.RST_BAR 0 0.187903f
c_1406 XDFSR12.CLKI_BAR 0 0.35929f
c_1413 XDFSR12.XML0.N1 0 0.0363245f
c_1421 XDFSR12.XML0.N2 0 0.123269f
c_1429 XDFSR12.XML0.N4 0 0.0453169f
c_1438 XDFSR12.XSL0.N1 0 0.12236f
c_1454 XDFSR12.CLKI 0 0.30462f
c_1464 XDFSR12.XSL0.N2 0 0.190162f
c_1474 XDFSR12.XSL0.N3 0 0.0472116f
c_1483 XDFSR11.N 0 0.157317f
c_1498 XDFSR11.RST_BAR 0 0.187903f
c_1515 XDFSR11.CLKI_BAR 0 0.35929f
c_1522 XDFSR11.XML0.N1 0 0.0363245f
c_1530 XDFSR11.XML0.N2 0 0.123269f
c_1538 XDFSR11.XML0.N4 0 0.0453169f
c_1547 XDFSR11.XSL0.N1 0 0.12236f
c_1563 XDFSR11.CLKI 0 0.30462f
c_1573 XDFSR11.XSL0.N2 0 0.190162f
c_1583 XDFSR11.XSL0.N3 0 0.0472116f
c_1592 XDFSR10.N 0 0.157317f
c_1607 XDFSR10.RST_BAR 0 0.187903f
c_1624 XDFSR10.CLKI_BAR 0 0.35929f
c_1631 XDFSR10.XML0.N1 0 0.0363245f
c_1639 XDFSR10.XML0.N2 0 0.123269f
c_1647 XDFSR10.XML0.N4 0 0.0453169f
c_1656 XDFSR10.XSL0.N1 0 0.12236f
c_1672 XDFSR10.CLKI 0 0.30462f
c_1682 XDFSR10.XSL0.N2 0 0.190162f
c_1692 XDFSR10.XSL0.N3 0 0.0472116f
c_1701 XDFSR9.N 0 0.157317f
c_1716 XDFSR9.RST_BAR 0 0.187903f
c_1733 XDFSR9.CLKI_BAR 0 0.35929f
c_1740 XDFSR9.XML0.N1 0 0.0363245f
c_1748 XDFSR9.XML0.N2 0 0.123269f
c_1756 XDFSR9.XML0.N4 0 0.0453169f
c_1765 XDFSR9.XSL0.N1 0 0.12236f
c_1781 XDFSR9.CLKI 0 0.30462f
c_1791 XDFSR9.XSL0.N2 0 0.190162f
c_1801 XDFSR9.XSL0.N3 0 0.0472116f
c_1810 XDFSR8.N 0 0.157317f
c_1825 XDFSR8.RST_BAR 0 0.187903f
c_1842 XDFSR8.CLKI_BAR 0 0.35929f
c_1849 XDFSR8.XML0.N1 0 0.0363245f
c_1857 XDFSR8.XML0.N2 0 0.123269f
c_1865 XDFSR8.XML0.N4 0 0.0453169f
c_1874 XDFSR8.XSL0.N1 0 0.12236f
c_1890 XDFSR8.CLKI 0 0.30462f
c_1900 XDFSR8.XSL0.N2 0 0.190162f
c_1910 XDFSR8.XSL0.N3 0 0.0472116f
c_1919 XDFSR7.N 0 0.157317f
c_1934 XDFSR7.RST_BAR 0 0.187903f
c_1951 XDFSR7.CLKI_BAR 0 0.35929f
c_1958 XDFSR7.XML0.N1 0 0.0363245f
c_1966 XDFSR7.XML0.N2 0 0.123269f
c_1974 XDFSR7.XML0.N4 0 0.0453169f
c_1983 XDFSR7.XSL0.N1 0 0.12236f
c_1999 XDFSR7.CLKI 0 0.30462f
c_2009 XDFSR7.XSL0.N2 0 0.190162f
c_2019 XDFSR7.XSL0.N3 0 0.0472116f
c_2028 XDFSR6.N 0 0.157317f
c_2043 XDFSR6.RST_BAR 0 0.187903f
c_2060 XDFSR6.CLKI_BAR 0 0.35929f
c_2067 XDFSR6.XML0.N1 0 0.0363245f
c_2075 XDFSR6.XML0.N2 0 0.123269f
c_2083 XDFSR6.XML0.N4 0 0.0453169f
c_2092 XDFSR6.XSL0.N1 0 0.12236f
c_2108 XDFSR6.CLKI 0 0.30462f
c_2118 XDFSR6.XSL0.N2 0 0.190162f
c_2128 XDFSR6.XSL0.N3 0 0.0472116f
c_2137 XDFSR5.N 0 0.157317f
c_2152 XDFSR5.RST_BAR 0 0.187159f
c_2169 XDFSR5.CLKI_BAR 0 0.35929f
c_2176 XDFSR5.XML0.N1 0 0.0363245f
c_2184 XDFSR5.XML0.N2 0 0.123269f
c_2192 XDFSR5.XML0.N4 0 0.0453169f
c_2201 XDFSR5.XSL0.N1 0 0.12236f
c_2217 XDFSR5.CLKI 0 0.30462f
c_2227 XDFSR5.XSL0.N2 0 0.190162f
c_2237 XDFSR5.XSL0.N3 0 0.0472116f
c_2247 XDFSR4.N 0 0.142219f
c_2263 XDFSR4.RST_BAR 0 0.159052f
c_2280 XDFSR4.CLKI_BAR 0 0.353979f
c_2287 XDFSR4.XML0.N1 0 0.0361574f
c_2296 XDFSR4.XML0.N2 0 0.120884f
c_2305 XDFSR4.XML0.N4 0 0.045049f
c_2315 XDFSR4.XSL0.N1 0 0.121163f
c_2331 XDFSR4.CLKI 0 0.295097f
c_2342 XDFSR4.XSL0.N2 0 0.189055f
c_2353 XDFSR4.XSL0.N3 0 0.0438555f
c_2363 XDFSR3.N 0 0.142219f
c_2379 XDFSR3.RST_BAR 0 0.159052f
c_2397 XDFSR3.CLKI_BAR 0 0.353979f
c_2405 XDFSR3.XML0.N1 0 0.0363245f
c_2414 XDFSR3.XML0.N2 0 0.121028f
c_2423 XDFSR3.XML0.N4 0 0.045049f
c_2433 XDFSR3.XSL0.N1 0 0.121163f
c_2450 XDFSR3.CLKI 0 0.295097f
c_2461 XDFSR3.XSL0.N2 0 0.189055f
c_2472 XDFSR3.XSL0.N3 0 0.0438555f
c_2483 XDFSR2.N 0 0.135695f
c_2500 XDFSR2.RST_BAR 0 0.154197f
c_2518 XDFSR2.CLKI_BAR 0 0.344763f
c_2526 XDFSR2.XML0.N1 0 0.0333679f
c_2536 XDFSR2.XML0.N2 0 0.118646f
c_2546 XDFSR2.XML0.N4 0 0.0434147f
c_2557 XDFSR2.XSL0.N1 0 0.118914f
c_2574 XDFSR2.CLKI 0 0.285757f
c_2586 XDFSR2.XSL0.N2 0 0.181953f
c_2598 XDFSR2.XSL0.N3 0 0.042543f
c_2610 XDFSR1.N 0 0.133503f
c_2628 XDFSR1.RST_BAR 0 0.151948f
c_2647 XDFSR1.CLKI_BAR 0 0.330538f
c_2656 XDFSR1.XML0.N1 0 0.0319055f
c_2667 XDFSR1.XML0.N2 0 0.116578f
c_2678 XDFSR1.XML0.N4 0 0.0429639f
c_2690 XDFSR1.XSL0.N1 0 0.116488f
c_2708 XDFSR1.CLKI 0 0.266575f
c_2721 XDFSR1.XSL0.N2 0 0.174505f
c_2734 XDFSR1.XSL0.N3 0 0.0433914f
c_2746 XDFSR0.N 0 0.133452f
c_2763 XDFSR0.RST_BAR 0 0.153594f
c_2783 XDFSR0.CLKI_BAR 0 0.332852f
c_2793 XDFSR0.XML0.N1 0 0.0319702f
c_2804 XDFSR0.XML0.N2 0 0.116711f
c_2815 XDFSR0.XML0.N4 0 0.0429444f
c_2827 XDFSR0.XSL0.N1 0 0.116488f
c_2845 XDFSR0.CLKI 0 0.268686f
c_2859 XDFSR0.XSL0.N2 0 0.171681f
c_2872 XDFSR0.XSL0.N3 0 0.0434508f
*
.include "LFSR.pex.netlist.LFSR.pxi"
*
.ends
*
*
