** Generated for: hspiceD
** Generated on: Dec  3 16:27:17 2021
** Design library name: cad6
** Design cell name: ALU_NO_FLAGS
** Design view name: schematic
.GLOBAL vdd! vss!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad6
** Cell name: NAND2_X1
** View name: schematic
.subckt NAND2_X1 a1 a2 zn
m_i_3 zn a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_2 vdd! a1 zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 zn a1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 net_0 a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends NAND2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: XNOR2_X1
** View name: schematic
.subckt XNOR2_X1 a b zn
m_i_48 net_003 a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_53 vdd! b net_003 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_29 net_000 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_36 vdd! b net_000 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_42 zn net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_0 net_001 a net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_5 vss! b net_001 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_11 net_002 net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_17 zn a net_002 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_23 net_002 b zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends XNOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: NOR2_X1
** View name: schematic
.subckt NOR2_X1 a1 a2 zn
m_i_1 zn a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 vss! a1 zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_2 zn a1 net_0 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_3 net_0 a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends NOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: MUX2_X1
** View name: schematic
.subckt MUX2_X1 a b s z
m_i_4 net_1 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_5 z_neg x1 net_1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_2 z_neg s net_0 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_3 net_0 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_10 vss! s x1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_6 net_2 s z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_8 vdd! a net_2 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_9 net_3 x1 z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_7 vdd! b net_3 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_11 vdd! s x1 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends MUX2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INV_X1
** View name: schematic
.subckt INV_X1 a zn
m_i_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: INVMUX2_X1
** View name: schematic
.subckt INVMUX2_X1 a b s zn
xi0 a b s z MUX2_X1
xi1 z zn INV_X1
.ends INVMUX2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: ALU_LOGIC_UNIT_1B
** View name: schematic
.subckt ALU_LOGIC_UNIT_1B ctrl<1> ctrl<0> logic_out op0 op1
xi0 op1 op0 nand_out NAND2_X1
xi1 op1 op0 xnor_out XNOR2_X1
xi2 op1 op0 nor_out NOR2_X1
xi4 nor_out op0 ctrl<0> mux1 MUX2_X1
xi3 nand_out xnor_out ctrl<0> mux0 MUX2_X1
xi5 mux0 mux1 ctrl<1> logic_out INVMUX2_X1
.ends ALU_LOGIC_UNIT_1B
** End of subcircuit definition.

** Library name: cad6
** Cell name: BUF_X1
** View name: schematic
.subckt BUF_X1 a z
m_i_3 vdd! a z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_2 vss! a z_neg vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends BUF_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: ALU_LOGIC_UNIT_16B
** View name: schematic
.subckt ALU_LOGIC_UNIT_16B ctrl<1> ctrl<0> logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> op0<15> op0<14> op0<13> op0<12> op0<11> op0<10> op0<9> op0<8> op0<7> op0<6> op0<5> op0<4> op0<3> op0<2> op0<1> op0<0> op1<15> op1<14> op1<13> op1<12> op1<11> op1<10> op1<9> op1<8> op1<7> op1<6> op1<5> op1<4> op1<3> op1<2> op1<1> op1<0>
xi18 ctrl1b<7> ctrl0b<7> logic_out<7> op0<7> op1<7> ALU_LOGIC_UNIT_1B
xi17 ctrl1b<3> ctrl0b<3> logic_out<3> op0<3> op1<3> ALU_LOGIC_UNIT_1B
xi16 ctrl1b<1> ctrl0b<1> logic_out<1> op0<1> op1<1> ALU_LOGIC_UNIT_1B
xi15 ctrl<1> ctrl<0> logic_out<0> op0<0> op1<0> ALU_LOGIC_UNIT_1B
xi14 ctrl1b<2> ctrl0b<2> logic_out<2> op0<2> op1<2> ALU_LOGIC_UNIT_1B
xi13 ctrl1b<5> ctrl0b<5> logic_out<5> op0<5> op1<5> ALU_LOGIC_UNIT_1B
xi0 ctrl1b<15> ctrl0b<15> logic_out<15> op0<15> op1<15> ALU_LOGIC_UNIT_1B
xi12 ctrl1b<4> ctrl0b<4> logic_out<4> op0<4> op1<4> ALU_LOGIC_UNIT_1B
xi11 ctrl1b<6> ctrl0b<6> logic_out<6> op0<6> op1<6> ALU_LOGIC_UNIT_1B
xi10 ctrl1b<11> ctrl0b<11> logic_out<11> op0<11> op1<11> ALU_LOGIC_UNIT_1B
xi9 ctrl1b<9> ctrl0b<9> logic_out<9> op0<9> op1<9> ALU_LOGIC_UNIT_1B
xi8 ctrl1b<8> ctrl0b<8> logic_out<8> op0<8> op1<8> ALU_LOGIC_UNIT_1B
xi7 ctrl1b<10> ctrl0b<10> logic_out<10> op0<10> op1<10> ALU_LOGIC_UNIT_1B
xi6 ctrl1b<13> ctrl0b<13> logic_out<13> op0<13> op1<13> ALU_LOGIC_UNIT_1B
xi5 ctrl1b<12> ctrl0b<12> logic_out<12> op0<12> op1<12> ALU_LOGIC_UNIT_1B
xi4 ctrl1b<14> ctrl0b<14> logic_out<14> op0<14> op1<14> ALU_LOGIC_UNIT_1B
xi33<1> ctrl1b<2> ctrl1b<3> BUF_X1
xi33<0> ctrl0b<2> ctrl0b<3> BUF_X1
xi32<1> ctrl1b<1> ctrl1b<2> BUF_X1
xi32<0> ctrl0b<1> ctrl0b<2> BUF_X1
xi31<1> ctrl<1> ctrl1b<1> BUF_X1
xi31<0> ctrl<0> ctrl0b<1> BUF_X1
xi30<1> ctrl1b<3> ctrl1b<4> BUF_X1
xi30<0> ctrl0b<3> ctrl0b<4> BUF_X1
xi24<1> ctrl1b<10> ctrl1b<11> BUF_X1
xi24<0> ctrl0b<10> ctrl0b<11> BUF_X1
xi23<1> ctrl1b<9> ctrl1b<10> BUF_X1
xi23<0> ctrl0b<9> ctrl0b<10> BUF_X1
xi22<1> ctrl1b<8> ctrl1b<9> BUF_X1
xi22<0> ctrl0b<8> ctrl0b<9> BUF_X1
xi29<1> ctrl1b<7> ctrl1b<8> BUF_X1
xi29<0> ctrl0b<7> ctrl0b<8> BUF_X1
xi28<1> ctrl1b<6> ctrl1b<7> BUF_X1
xi28<0> ctrl0b<6> ctrl0b<7> BUF_X1
xi27<1> ctrl1b<5> ctrl1b<6> BUF_X1
xi27<0> ctrl0b<5> ctrl0b<6> BUF_X1
xi26<1> ctrl1b<4> ctrl1b<5> BUF_X1
xi26<0> ctrl0b<4> ctrl0b<5> BUF_X1
xi25<1> ctrl1b<11> ctrl1b<12> BUF_X1
xi25<0> ctrl0b<11> ctrl0b<12> BUF_X1
xi19<1> ctrl1b<14> ctrl1b<15> BUF_X1
xi19<0> ctrl0b<14> ctrl0b<15> BUF_X1
xi21<1> ctrl1b<13> ctrl1b<14> BUF_X1
xi21<0> ctrl0b<13> ctrl0b<14> BUF_X1
xi20<1> ctrl1b<12> ctrl1b<13> BUF_X1
xi20<0> ctrl0b<12> ctrl0b<13> BUF_X1
.ends ALU_LOGIC_UNIT_16B
** End of subcircuit definition.

** Library name: cad6
** Cell name: FA_X1
** View name: schematic
.subckt FA_X1 a b ci co s
m_instance_284 net_010 ci net_005 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_280 net_009 b net_010 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_275 vdd! a net_009 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_251 net_007 a net_001 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_246 vdd! b net_007 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_239 co net_001 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_instance_315 s net_005 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_269 net_008 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_263 vdd! b net_008 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_257 net_001 ci net_008 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_309 net_011 b vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_297 vdd! ci net_011 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_303 net_011 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_290 net_005 net_001 net_011 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_203 net_004 ci net_005 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_199 net_003 b net_004 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_194 vss! a net_003 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_159 co net_001 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_233 s net_005 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_166 vss! b net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_170 net_000 a net_001 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_176 net_001 ci net_002 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_209 net_005 net_001 net_006 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_215 vss! ci net_006 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_188 net_002 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_182 vss! b net_002 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_227 net_006 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_221 net_006 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
.ends FA_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: XOR2_X1
** View name: schematic
.subckt XOR2_X1 a b z
m_i_19 net_001 a z vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_24 vss! b net_001 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0 net_000 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_13 z net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_7 vss! b net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_30 net_002 a net_000 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_35 vdd! b net_002 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_41 net_003 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_47 z a net_003 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_53 net_003 b z vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends XOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: RCA_4B
** View name: schematic
.subckt RCA_4B co logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> s<3> s<2> s<1> s<0> ctrl<0> ctrl_out<0> op0<3> op0<2> op0<1> op0<0> op1<3> op1<2> op1<1> op1<0>
xi3 op0_temp<3> op1<3> net26 net1 s<3> FA_X1
xi2 op0_temp<2> op1<2> net21 net26 s<2> FA_X1
xi1 op0_temp<1> op1<1> net16 net21 s<1> FA_X1
xi0 op0_temp<0> op1<0> ctrl<0> net16 s<0> FA_X1
xi12 ctrl_buf<3> op0<3> op0_temp<3> XOR2_X1
xi11 ctrl_buf<2> op0<2> op0_temp<2> XOR2_X1
xi10 ctrl_buf<1> op0<1> op0_temp<1> XOR2_X1
xi9 ctrl<0> op0<0> op0_temp<0> XOR2_X1
xi29 net1 co BUF_X1
xi19<3> logic_out<3> logic_out_buf<3> BUF_X1
xi19<2> logic_out<2> logic_out_buf<2> BUF_X1
xi19<1> logic_out<1> logic_out_buf<1> BUF_X1
xi19<0> logic_out<0> logic_out_buf<0> BUF_X1
xi16 ctrl_buf<2> ctrl_buf<3> BUF_X1
xi15 ctrl_buf<1> ctrl_buf<2> BUF_X1
xi14 ctrl<0> ctrl_buf<1> BUF_X1
xi13 ctrl_buf<3> ctrl_out<0> BUF_X1
.ends RCA_4B
** End of subcircuit definition.

** Library name: cad6
** Cell name: CSA_4B
** View name: schematic
.subckt CSA_4B ci co logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> s<3> s<2> s<1> s<0> ctrl<0> ctrl_out<0> op0<3> op0<2> op0<1> op0<0> op0_temp<3> op1<3> op1<2> op1<1> op1<0>
xi8 op0_temp<3> op1<3> net46 co_1 s_1<3> FA_X1
xi7 op0_temp<2> op1<2> net41 net46 s_1<2> FA_X1
xi6 op0_temp<1> op1<1> net36 net41 s_1<1> FA_X1
xi5 op0_temp<0> op1<0> vdd! net36 s_1<0> FA_X1
xi3 op0_temp<3> op1<3> net26 co_0 s_0<3> FA_X1
xi2 op0_temp<2> op1<2> net21 net26 s_0<2> FA_X1
xi1 op0_temp<1> op1<1> net16 net21 s_0<1> FA_X1
xi0 op0_temp<0> op1<0> vss! net16 s_0<0> FA_X1
xi12 ctrl_buf<3> op0<3> op0_temp<3> XOR2_X1
xi11 ctrl_buf<2> op0<2> op0_temp<2> XOR2_X1
xi10 ctrl_buf<1> op0<1> op0_temp<1> XOR2_X1
xi9 ctrl<0> op0<0> op0_temp<0> XOR2_X1
xi28 ci_buf<3> ci_buf_s_co BUF_X1
xi21 ci ci_buf<1> BUF_X1
xi19<3> logic_out<3> logic_out_buf<3> BUF_X1
xi19<2> logic_out<2> logic_out_buf<2> BUF_X1
xi19<1> logic_out<1> logic_out_buf<1> BUF_X1
xi19<0> logic_out<0> logic_out_buf<0> BUF_X1
xi20 ci_buf<1> ci_buf<2> BUF_X1
xi27 ci_buf<2> ci_buf<3> BUF_X1
xi16 ctrl_buf<2> ctrl_buf<3> BUF_X1
xi15 ctrl_buf<1> ctrl_buf<2> BUF_X1
xi14 ctrl<0> ctrl_buf<1> BUF_X1
xi13 ctrl_buf<3> ctrl_out<0> BUF_X1
xi17 s_0<0> s_1<0> ci s<0> MUX2_X1
xi24 s_0<3> s_1<3> ci_buf<3> s<3> MUX2_X1
xi26 s_0<2> s_1<2> ci_buf<2> s<2> MUX2_X1
xi25 s_0<1> s_1<1> ci_buf<1> s<1> MUX2_X1
xi18 co_0 co_1 ci_buf_s_co co MUX2_X1
.ends CSA_4B
** End of subcircuit definition.

** Library name: cad6
** Cell name: ALU_ARITHMETIC_UNIT_16B
** View name: schematic
.subckt ALU_ARITHMETIC_UNIT_16B arithmetic_out<15> arithmetic_out<14> arithmetic_out<13> arithmetic_out<12> arithmetic_out<11> arithmetic_out<10> arithmetic_out<9> arithmetic_out<8> arithmetic_out<7> arithmetic_out<6> arithmetic_out<5> arithmetic_out<4> arithmetic_out<3> arithmetic_out<2> arithmetic_out<1> arithmetic_out<0> co logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<15> logic_out_buf<14> logic_out_buf<13> logic_out_buf<12> logic_out_buf<11> logic_out_buf<10> logic_out_buf<9> logic_out_buf<8> logic_out_buf<7> logic_out_buf<6> logic_out_buf<5> logic_out_buf<4> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> ctrl<0> op0<15> op0<14> op0<13> op0<12> op0<11> op0<10> op0<9> op0<8> op0<7> op0<6> op0<5> op0<4> op0<3> op0<2> op0<1> op0<0> op0_temp<15> op1<15> op1<14> op1<13> op1<12> op1<11> op1<10> op1<9> op1<8>
+op1<7> op1<6> op1<5> op1<4> op1<3> op1<2> op1<1> op1<0>
xi3 net1 logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> arithmetic_out<3> arithmetic_out<2> arithmetic_out<1> arithmetic_out<0> ctrl<0> net3 op0<3> op0<2> op0<1> op0<0> op1<3> op1<2> op1<1> op1<0> RCA_4B
xi4 net1 net4 logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out_buf<7> logic_out_buf<6> logic_out_buf<5> logic_out_buf<4> arithmetic_out<7> arithmetic_out<6> arithmetic_out<5> arithmetic_out<4> net3 net7 op0<7> op0<6> op0<5> op0<4> net10 op1<7> op1<6> op1<5> op1<4> CSA_4B
xi6 net5 co logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out_buf<15> logic_out_buf<14> logic_out_buf<13> logic_out_buf<12> arithmetic_out<15> arithmetic_out<14> arithmetic_out<13> arithmetic_out<12> net8 net9 op0<15> op0<14> op0<13> op0<12> op0_temp<15> op1<15> op1<14> op1<13> op1<12> CSA_4B
xi5 net4 net5 logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out_buf<11> logic_out_buf<10> logic_out_buf<9> logic_out_buf<8> arithmetic_out<11> arithmetic_out<10> arithmetic_out<9> arithmetic_out<8> net7 net8 op0<11> op0<10> op0<9> op0<8> net6 op1<11> op1<10> op1<9> op1<8> CSA_4B
.ends ALU_ARITHMETIC_UNIT_16B
** End of subcircuit definition.

** Library name: cad6
** Cell name: INV_X4
** View name: schematic
.subckt INV_X4 a zn
m_i_1_0_x4_0 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_1 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_2 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_1_0_x4_3 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0_0_x4_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_1 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_2 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0_0_x4_3 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV_X4
** End of subcircuit definition.

** Library name: cad6
** Cell name: OUT_MUX_BUF_16B
** View name: schematic
.subckt OUT_MUX_BUF_16B arithmetic_out<15> arithmetic_out<14> arithmetic_out<13> arithmetic_out<12> arithmetic_out<11> arithmetic_out<10> arithmetic_out<9> arithmetic_out<8> arithmetic_out<7> arithmetic_out<6> arithmetic_out<5> arithmetic_out<4> arithmetic_out<3> arithmetic_out<2> arithmetic_out<1> arithmetic_out<0> logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> alu_out<15> alu_out<14> alu_out<13> alu_out<12> alu_out<11> alu_out<10> alu_out<9> alu_out<8> alu_out<7> alu_out<6> alu_out<5> alu_out<4> alu_out<3> alu_out<2> alu_out<1> alu_out<0> alu_pre<15> ctrl<2>
xi0<15> logic_out<15> arithmetic_out<15> ctrl_2_buf<15> alu_pre<15> MUX2_X1
xi0<14> logic_out<14> arithmetic_out<14> ctrl_2_buf<14> alu_pre<14> MUX2_X1
xi0<13> logic_out<13> arithmetic_out<13> ctrl_2_buf<13> alu_pre<13> MUX2_X1
xi0<12> logic_out<12> arithmetic_out<12> ctrl_2_buf<12> alu_pre<12> MUX2_X1
xi0<11> logic_out<11> arithmetic_out<11> ctrl_2_buf<11> alu_pre<11> MUX2_X1
xi0<10> logic_out<10> arithmetic_out<10> ctrl_2_buf<10> alu_pre<10> MUX2_X1
xi0<9> logic_out<9> arithmetic_out<9> ctrl_2_buf<9> alu_pre<9> MUX2_X1
xi0<8> logic_out<8> arithmetic_out<8> ctrl_2_buf<8> alu_pre<8> MUX2_X1
xi0<7> logic_out<7> arithmetic_out<7> ctrl_2_buf<7> alu_pre<7> MUX2_X1
xi0<6> logic_out<6> arithmetic_out<6> ctrl_2_buf<6> alu_pre<6> MUX2_X1
xi0<5> logic_out<5> arithmetic_out<5> ctrl_2_buf<5> alu_pre<5> MUX2_X1
xi0<4> logic_out<4> arithmetic_out<4> ctrl_2_buf<4> alu_pre<4> MUX2_X1
xi0<3> logic_out<3> arithmetic_out<3> ctrl_2_buf<3> alu_pre<3> MUX2_X1
xi0<2> logic_out<2> arithmetic_out<2> ctrl_2_buf<2> alu_pre<2> MUX2_X1
xi0<1> logic_out<1> arithmetic_out<1> ctrl_2_buf<1> alu_pre<1> MUX2_X1
xi0<0> logic_out<0> arithmetic_out<0> ctrl_2_buf<0> alu_pre<0> MUX2_X1
xi1<15> alu_pre<15> net3<0> INV_X1
xi1<14> alu_pre<14> net3<1> INV_X1
xi1<13> alu_pre<13> net3<2> INV_X1
xi1<12> alu_pre<12> net3<3> INV_X1
xi1<11> alu_pre<11> net3<4> INV_X1
xi1<10> alu_pre<10> net3<5> INV_X1
xi1<9> alu_pre<9> net3<6> INV_X1
xi1<8> alu_pre<8> net3<7> INV_X1
xi1<7> alu_pre<7> net3<8> INV_X1
xi1<6> alu_pre<6> net3<9> INV_X1
xi1<5> alu_pre<5> net3<10> INV_X1
xi1<4> alu_pre<4> net3<11> INV_X1
xi1<3> alu_pre<3> net3<12> INV_X1
xi1<2> alu_pre<2> net3<13> INV_X1
xi1<1> alu_pre<1> net3<14> INV_X1
xi1<0> alu_pre<0> net3<15> INV_X1
xi2<15> net3<0> alu_out<15> INV_X4
xi2<14> net3<1> alu_out<14> INV_X4
xi2<13> net3<2> alu_out<13> INV_X4
xi2<12> net3<3> alu_out<12> INV_X4
xi2<11> net3<4> alu_out<11> INV_X4
xi2<10> net3<5> alu_out<10> INV_X4
xi2<9> net3<6> alu_out<9> INV_X4
xi2<8> net3<7> alu_out<8> INV_X4
xi2<7> net3<8> alu_out<7> INV_X4
xi2<6> net3<9> alu_out<6> INV_X4
xi2<5> net3<10> alu_out<5> INV_X4
xi2<4> net3<11> alu_out<4> INV_X4
xi2<3> net3<12> alu_out<3> INV_X4
xi2<2> net3<13> alu_out<2> INV_X4
xi2<1> net3<14> alu_out<1> INV_X4
xi2<0> net3<15> alu_out<0> INV_X4
xi27 ctrl_2_buf<13> ctrl_2_buf<12> BUF_X1
xi26 ctrl_2_buf<14> ctrl_2_buf<13> BUF_X1
xi25 ctrl_2_buf<15> ctrl_2_buf<14> BUF_X1
xi24 ctrl<2> ctrl_2_buf<15> BUF_X1
xi23 ctrl_2_buf<12> ctrl_2_buf<11> BUF_X1
xi22 ctrl_2_buf<11> ctrl_2_buf<10> BUF_X1
xi21 ctrl_2_buf<10> ctrl_2_buf<9> BUF_X1
xi20 ctrl_2_buf<9> ctrl_2_buf<8> BUF_X1
xi19 ctrl_2_buf<5> ctrl_2_buf<4> BUF_X1
xi18 ctrl_2_buf<6> ctrl_2_buf<5> BUF_X1
xi17 ctrl_2_buf<7> ctrl_2_buf<6> BUF_X1
xi16 ctrl_2_buf<8> ctrl_2_buf<7> BUF_X1
xi12 ctrl_2_buf<4> ctrl_2_buf<3> BUF_X1
xi11 ctrl_2_buf<3> ctrl_2_buf<2> BUF_X1
xi4 ctrl_2_buf<2> ctrl_2_buf<1> BUF_X1
xi3 ctrl_2_buf<1> ctrl_2_buf<0> BUF_X1
.ends OUT_MUX_BUF_16B
** End of subcircuit definition.

** Library name: cad6
** Cell name: ALU_NO_FLAGS
** View name: schematic
xi0 ctrl<1> ctrl<0> logic_pre<15> logic_pre<14> logic_pre<13> logic_pre<12> logic_pre<11> logic_pre<10> logic_pre<9> logic_pre<8> logic_pre<7> logic_pre<6> logic_pre<5> logic_pre<4> logic_pre<3> logic_pre<2> logic_pre<1> logic_pre<0> op0<15> op0<14> op0<13> op0<12> op0<11> op0<10> op0<9> op0<8> op0<7> op0<6> op0<5> op0<4> op0<3> op0<2> op0<1> op0<0> op1<15> op1<14> op1<13> op1<12> op1<11> op1<10> op1<9> op1<8> op1<7> op1<6> op1<5> op1<4> op1<3> op1<2> op1<1> op1<0> ALU_LOGIC_UNIT_16B
xi1 arithmetic_out<15> arithmetic_out<14> arithmetic_out<13> arithmetic_out<12> arithmetic_out<11> arithmetic_out<10> arithmetic_out<9> arithmetic_out<8> arithmetic_out<7> arithmetic_out<6> arithmetic_out<5> arithmetic_out<4> arithmetic_out<3> arithmetic_out<2> arithmetic_out<1> arithmetic_out<0> co logic_pre<15> logic_pre<14> logic_pre<13> logic_pre<12> logic_pre<11> logic_pre<10> logic_pre<9> logic_pre<8> logic_pre<7> logic_pre<6> logic_pre<5> logic_pre<4> logic_pre<3> logic_pre<2> logic_pre<1> logic_pre<0> logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> ctrl<0> op0<15> op0<14> op0<13> op0<12> op0<11> op0<10> op0<9> op0<8> op0<7> op0<6> op0<5> op0<4> op0<3> op0<2> op0<1> op0<0> op0_temp<15> op1<15> op1<14> op1<13> op1<12> op1<11> op1<10> op1<9> op1<8> op1<7> op1<6> op1<5> op1<4> op1<3> op1<2> op1<1> op1<0> ALU_ARITHMETIC_UNIT_16B
xi2 arithmetic_out<15> arithmetic_out<14> arithmetic_out<13> arithmetic_out<12> arithmetic_out<11> arithmetic_out<10> arithmetic_out<9> arithmetic_out<8> arithmetic_out<7> arithmetic_out<6> arithmetic_out<5> arithmetic_out<4> arithmetic_out<3> arithmetic_out<2> arithmetic_out<1> arithmetic_out<0> logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out<3> logic_out<2> logic_out<1> logic_out<0> alu_out<15> alu_out<14> alu_out<13> alu_out<12> alu_out<11> alu_out<10> alu_out<9> alu_out<8> alu_out<7> alu_out<6> alu_out<5> alu_out<4> alu_out<3> alu_out<2> alu_out<1> alu_out<0> alu_pre<15> ctrl<2> OUT_MUX_BUF_16B
.END
