
* Subcircuits
*---------------------------------------------------------------------------------------------------
.INCLUDE 'INV1.ckt'
*---------------------------------------------------------------------------------------------------
.subckt BUF1 in out vdd vss M=1
xi0 in n1 vdd vss INV1 
xi1 n1 out vdd vss INV1 
.ends BUF1
