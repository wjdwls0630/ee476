../../netlist/PEX/penalty.pex.netlist