** Generated for: hspiceD
** Generated on: Nov 12 21:24:22 2021
** Design library name: cad5
** Design cell name: T2BREG_LATCH
** Design view name: schematic
.GLOBAL vss! vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad5
** Cell name: INV_X4
** View name: schematic
.subckt INV_X4 a zn
m_i_0_0_x4_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_0_x4_1 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_0_x4_2 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_0_x4_3 vss! a zn vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1_0_x4_0 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_1_0_x4_1 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_1_0_x4_2 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_1_0_x4_3 vdd! a zn vdd! PMOS_VTL L=50e-9 W=630e-9
.ends INV_X4
** End of subcircuit definition.

** Library name: cad5
** Cell name: INV_X1
** View name: schematic
.subckt INV_X1 a zn
m_i_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
.ends INV_X1
** End of subcircuit definition.

** Library name: cad5
** Cell name: DLL_X1
** View name: schematic
.subckt DLL_X1 d gn q
m_i_13 net_002 d vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_18 net_003 net_000 net_002 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_24 net_004 net_001 net_003 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_29 vss! net_005 net_004 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_42 q net_003 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0 net_000 gn vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_7 vss! net_000 net_001 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_35 vss! net_003 net_005 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_67 net_003 net_001 net_006 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_62 net_006 d vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_79 vdd! net_005 net_007 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_73 net_007 net_000 net_003 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_92 q net_003 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_48 net_000 gn vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_55 vdd! net_000 net_001 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_85 vdd! net_003 net_005 vdd! PMOS_VTL L=50e-9 W=90e-9
.ends DLL_X1
** End of subcircuit definition.

** Library name: cad5
** Cell name: TBUF_X2
** View name: schematic
.subckt TBUF_X2 a en z
m_i_0_15_63 dummy1 a y vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_14_47 vss! nen dummy1 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_15 vss! a x vss! NMOS_VTL L=50e-9 W=415e-9
m_i_17 vss! en nen vss! NMOS_VTL L=50e-9 W=210e-9
m_i_0_14 vss! en x vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0_6 vss! x z vss! NMOS_VTL L=50e-9 W=355e-9
m_i_0 vss! x z vss! NMOS_VTL L=50e-9 W=355e-9
m_i_24_1 dummy0 en x vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_24_0 vdd! a dummy0 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_24_0_64 vdd! a y vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_24_3 vdd! y z vdd! PMOS_VTL L=50e-9 W=540e-9
m_i_24 vdd! y z vdd! PMOS_VTL L=50e-9 W=540e-9
m_i_24_1_48 y nen vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_42 vdd! en nen vdd! PMOS_VTL L=50e-9 W=315e-9
.ends TBUF_X2
** End of subcircuit definition.

** Library name: cad5
** Cell name: DLH_X1
** View name: schematic
.subckt DLH_X1 d g q
m_i_13 net_002 d vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_18 net_003 net_001 net_002 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_28 vss! net_005 net_004 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_24 net_004 net_000 net_003 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_0 vss! g net_000 vss! NMOS_VTL L=50e-9 W=210e-9
m_i_41_11 q net_003 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_7 net_001 net_000 vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_i_34 vss! net_003 net_005 vss! NMOS_VTL L=50e-9 W=90e-9
m_i_66 net_003 net_000 net_006 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_61 net_006 d vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_72 net_007 net_001 net_003 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_76 vdd! net_005 net_007 vdd! PMOS_VTL L=50e-9 W=90e-9
m_i_48 vdd! g net_000 vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_89_4 q net_003 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_55 net_001 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_i_82 vdd! net_003 net_005 vdd! PMOS_VTL L=50e-9 W=90e-9
.ends DLH_X1
** End of subcircuit definition.

** Library name: cad5
** Cell name: T2BREG_LATCH
** View name: schematic
xi12<1> wr_data_preinv<1> wr_data_b<1> INV_X4
xi12<0> wr_data_preinv<0> wr_data_b<0> INV_X4
xi11<1> wr_data_prebuff<1> wr_data_preinv<1> INV_X1
xi11<0> wr_data_prebuff<0> wr_data_preinv<0> INV_X1
xi6<1> wr_data<1> ck wr_data_prebuff<1> DLL_X1
xi6<0> wr_data<0> ck wr_data_prebuff<0> DLL_X1
xi10<1> reg_data_1<1> r1_d1 rd_data_1<1> TBUF_X2
xi10<0> reg_data_1<0> r1_d1 rd_data_1<0> TBUF_X2
xi9<1> reg_data_1<1> r0_d1 rd_data_0<1> TBUF_X2
xi9<0> reg_data_1<0> r0_d1 rd_data_0<0> TBUF_X2
xi3<1> reg_data_0<1> r1_d0 rd_data_1<1> TBUF_X2
xi3<0> reg_data_0<0> r1_d0 rd_data_1<0> TBUF_X2
xi4<1> reg_data_0<1> r0_d0 rd_data_0<1> TBUF_X2
xi4<0> reg_data_0<0> r0_d0 rd_data_0<0> TBUF_X2
xi8<1> wr_data_b<1> ck_1 reg_data_1<1> DLH_X1
xi8<0> wr_data_b<0> ck_1 reg_data_1<0> DLH_X1
xi7<1> wr_data_b<1> ck_0 reg_data_0<1> DLH_X1
xi7<0> wr_data_b<0> ck_0 reg_data_0<0> DLH_X1
.END
