* File: ring_osc.pex.netlist
* Created: Fri Oct 29 05:27:39 2021
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.subckt ring_osc_pex OSC_EN OSC_OUT
* 
mXI0.MNMOS0 XI0.NET2 OSC_EN VSS! VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI0.MNMOS1 NET3 OSC_OUT XI0.NET2 VSS! NMOS_VTG L=6e-08 W=3.5e-07 AD=3.675e-14
+ AS=5.6e-14 PD=9.1e-07 PS=1.02e-06
mXI0.MPMOS0 NET3 OSC_EN VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI0.MPMOS1 NET3 OSC_OUT VDD! VDD! PMOS_VTG L=6e-08 W=3.5e-07 AD=5.6e-14
+ AS=3.675e-14 PD=1.02e-06 PS=9.1e-07
mXI8.MM0 OSC_OUT NET17 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14
+ AS=3.15e-14 PD=8.1e-07 PS=8.1e-07
mXI8.MM1 OSC_OUT NET17 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI1.MM0 NET5 NET3 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI1.MM1 NET5 NET3 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI7.MM0 NET17 NET15 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI7.MM1 NET17 NET15 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI2.MM0 NET7 NET5 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI2.MM1 NET7 NET5 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI6.MM0 NET15 NET13 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI6.MM1 NET15 NET13 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI3.MM0 NET9 NET7 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI3.MM1 NET9 NET7 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI5.MM0 NET13 NET11 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI5.MM1 NET13 NET11 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
mXI4.MM0 NET11 NET9 VSS! VSS! NMOS_VTG L=6e-08 W=3e-07 AD=3.15e-14 AS=3.15e-14
+ PD=8.1e-07 PS=8.1e-07
mXI4.MM1 NET11 NET9 VDD! VDD! PMOS_VTG L=6e-08 W=4e-07 AD=4.2e-14 AS=4.2e-14
+ PD=1.01e-06 PS=1.01e-06
c_7 OSC_OUT 0 0.161923f
c_19 VDD! 0 0.487277f
c_24 NET11 0 0.201042f
c_29 OSC_EN 0 0.0666759f
c_41 VSS! 0 0.177173f
c_47 NET3 0 0.130375f
c_52 NET17 0 0.0983505f
c_58 NET5 0 0.0984607f
c_63 NET15 0 0.0881648f
c_68 NET7 0 0.0844663f
c_73 NET13 0 0.0926826f
c_78 NET9 0 0.0947361f
*
.include "ring_osc.pex.netlist.RING_OSC.pxi"
*
.ends
*
*
