** Generated for: hspiceD
** Generated on: Dec  3 16:28:11 2021
** Design library name: cad6
** Design cell name: ALU_ARITHMETIC_UNIT_16B
** Design view name: schematic
.GLOBAL vss! vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad6
** Cell name: FA_X1
** View name: schematic
.subckt FA_X1 a b ci co s
m_instance_284 net_010 ci net_005 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_280 net_009 b net_010 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_275 vdd! a net_009 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_251 net_007 a net_001 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_246 vdd! b net_007 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_239 co net_001 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_instance_315 s net_005 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_269 net_008 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_263 vdd! b net_008 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_257 net_001 ci net_008 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_309 net_011 b vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_297 vdd! ci net_011 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_303 net_011 a vdd! vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_290 net_005 net_001 net_011 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_instance_203 net_004 ci net_005 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_199 net_003 b net_004 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_194 vss! a net_003 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_159 co net_001 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_233 s net_005 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_166 vss! b net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_170 net_000 a net_001 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_176 net_001 ci net_002 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_209 net_005 net_001 net_006 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_215 vss! ci net_006 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_188 net_002 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_182 vss! b net_002 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_instance_227 net_006 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_instance_221 net_006 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
.ends FA_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: XOR2_X1
** View name: schematic
.subckt XOR2_X1 a b z
m_i_19 net_001 a z vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_24 vss! b net_001 vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_0 net_000 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_13 z net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=43.575e-15 AS=43.575e-15 PD=625e-9 PS=625e-9 M=1
m_i_7 vss! b net_000 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_30 net_002 a net_000 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_35 vdd! b net_002 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_41 net_003 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=66.15e-15 AS=66.15e-15 PD=840e-9 PS=840e-9 M=1
m_i_47 z a net_003 vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_53 net_003 b z vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends XOR2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: BUF_X1
** View name: schematic
.subckt BUF_X1 a z
m_i_3 vdd! a z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_2 vss! a z_neg vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends BUF_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: RCA_4B
** View name: schematic
.subckt RCA_4B co logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> s<3> s<2> s<1> s<0> ctrl<0> ctrl_out<0> op0<3> op0<2> op0<1> op0<0> op1<3> op1<2> op1<1> op1<0>
xi3 op0_temp<3> op1<3> net26 net1 s<3> FA_X1
xi2 op0_temp<2> op1<2> net21 net26 s<2> FA_X1
xi1 op0_temp<1> op1<1> net16 net21 s<1> FA_X1
xi0 op0_temp<0> op1<0> ctrl<0> net16 s<0> FA_X1
xi12 ctrl_buf<3> op0<3> op0_temp<3> XOR2_X1
xi11 ctrl_buf<2> op0<2> op0_temp<2> XOR2_X1
xi10 ctrl_buf<1> op0<1> op0_temp<1> XOR2_X1
xi9 ctrl<0> op0<0> op0_temp<0> XOR2_X1
xi29 net1 co BUF_X1
xi19<3> logic_out<3> logic_out_buf<3> BUF_X1
xi19<2> logic_out<2> logic_out_buf<2> BUF_X1
xi19<1> logic_out<1> logic_out_buf<1> BUF_X1
xi19<0> logic_out<0> logic_out_buf<0> BUF_X1
xi16 ctrl_buf<2> ctrl_buf<3> BUF_X1
xi15 ctrl_buf<1> ctrl_buf<2> BUF_X1
xi14 ctrl<0> ctrl_buf<1> BUF_X1
xi13 ctrl_buf<3> ctrl_out<0> BUF_X1
.ends RCA_4B
** End of subcircuit definition.

** Library name: cad6
** Cell name: MUX2_X1
** View name: schematic
.subckt MUX2_X1 a b s z
m_i_4 net_1 a vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_5 z_neg x1 net_1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_2 z_neg s net_0 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_3 net_0 b vss! vss! NMOS_VTL L=50e-9 W=210e-9 AD=22.05e-15 AS=22.05e-15 PD=420e-9 PS=420e-9 M=1
m_i_0 z z_neg vss! vss! NMOS_VTL L=50e-9 W=415e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_10 vss! s x1 vss! NMOS_VTL L=50e-9 W=210e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_6 net_2 s z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_8 vdd! a net_2 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_9 net_3 x1 z_neg vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_7 vdd! b net_3 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=33.075e-15 AS=33.075e-15 PD=525e-9 PS=525e-9 M=1
m_i_1 z z_neg vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m_i_11 vdd! s x1 vdd! PMOS_VTL L=50e-9 W=315e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends MUX2_X1
** End of subcircuit definition.

** Library name: cad6
** Cell name: CSA_4B
** View name: schematic
.subckt CSA_4B ci co logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> s<3> s<2> s<1> s<0> ctrl<0> ctrl_out<0> op0<3> op0<2> op0<1> op0<0> op0_temp<3> op1<3> op1<2> op1<1> op1<0>
xi8 op0_temp<3> op1<3> net46 co_1 s_1<3> FA_X1
xi7 op0_temp<2> op1<2> net41 net46 s_1<2> FA_X1
xi6 op0_temp<1> op1<1> net36 net41 s_1<1> FA_X1
xi5 op0_temp<0> op1<0> vdd! net36 s_1<0> FA_X1
xi3 op0_temp<3> op1<3> net26 co_0 s_0<3> FA_X1
xi2 op0_temp<2> op1<2> net21 net26 s_0<2> FA_X1
xi1 op0_temp<1> op1<1> net16 net21 s_0<1> FA_X1
xi0 op0_temp<0> op1<0> vss! net16 s_0<0> FA_X1
xi12 ctrl_buf<3> op0<3> op0_temp<3> XOR2_X1
xi11 ctrl_buf<2> op0<2> op0_temp<2> XOR2_X1
xi10 ctrl_buf<1> op0<1> op0_temp<1> XOR2_X1
xi9 ctrl<0> op0<0> op0_temp<0> XOR2_X1
xi28 ci_buf<3> ci_buf_s_co BUF_X1
xi21 ci ci_buf<1> BUF_X1
xi19<3> logic_out<3> logic_out_buf<3> BUF_X1
xi19<2> logic_out<2> logic_out_buf<2> BUF_X1
xi19<1> logic_out<1> logic_out_buf<1> BUF_X1
xi19<0> logic_out<0> logic_out_buf<0> BUF_X1
xi20 ci_buf<1> ci_buf<2> BUF_X1
xi27 ci_buf<2> ci_buf<3> BUF_X1
xi16 ctrl_buf<2> ctrl_buf<3> BUF_X1
xi15 ctrl_buf<1> ctrl_buf<2> BUF_X1
xi14 ctrl<0> ctrl_buf<1> BUF_X1
xi13 ctrl_buf<3> ctrl_out<0> BUF_X1
xi17 s_0<0> s_1<0> ci s<0> MUX2_X1
xi24 s_0<3> s_1<3> ci_buf<3> s<3> MUX2_X1
xi26 s_0<2> s_1<2> ci_buf<2> s<2> MUX2_X1
xi25 s_0<1> s_1<1> ci_buf<1> s<1> MUX2_X1
xi18 co_0 co_1 ci_buf_s_co co MUX2_X1
.ends CSA_4B
** End of subcircuit definition.

** Library name: cad6
** Cell name: ALU_ARITHMETIC_UNIT_16B
** View name: schematic
xi3 net1 logic_out<3> logic_out<2> logic_out<1> logic_out<0> logic_out_buf<3> logic_out_buf<2> logic_out_buf<1> logic_out_buf<0> arithmetic_out<3> arithmetic_out<2> arithmetic_out<1> arithmetic_out<0> ctrl<0> net3 op0<3> op0<2> op0<1> op0<0> op1<3> op1<2> op1<1> op1<0> RCA_4B
xi4 net1 net4 logic_out<7> logic_out<6> logic_out<5> logic_out<4> logic_out_buf<7> logic_out_buf<6> logic_out_buf<5> logic_out_buf<4> arithmetic_out<7> arithmetic_out<6> arithmetic_out<5> arithmetic_out<4> net3 net7 op0<7> op0<6> op0<5> op0<4> net10 op1<7> op1<6> op1<5> op1<4> CSA_4B
xi6 net5 co logic_out<15> logic_out<14> logic_out<13> logic_out<12> logic_out_buf<15> logic_out_buf<14> logic_out_buf<13> logic_out_buf<12> arithmetic_out<15> arithmetic_out<14> arithmetic_out<13> arithmetic_out<12> net8 net9 op0<15> op0<14> op0<13> op0<12> op0_temp<15> op1<15> op1<14> op1<13> op1<12> CSA_4B
xi5 net4 net5 logic_out<11> logic_out<10> logic_out<9> logic_out<8> logic_out_buf<11> logic_out_buf<10> logic_out_buf<9> logic_out_buf<8> arithmetic_out<11> arithmetic_out<10> arithmetic_out<9> arithmetic_out<8> net7 net8 op0<11> op0<10> op0<9> op0<8> net6 op1<11> op1<10> op1<9> op1<8> CSA_4B
.END
