* 1   2   3   4
* in out en en_bar
.subckt TG_DFSR 1 2 3 4 Wp=0.4e-6 Wn=0.3e-6
mn0 1 3 2 vss! NMOS_VTG L=60e-9 W='Wn' AD='0.105e-6*Wn' AS='0.105e-6*Wn' PD='Wn+210e-9' PS='Wn+210e-9' M=1
mp0 1 4 2 vdd! PMOS_VTG L=60e-9 W='Wp' AD='0.105e-6*Wp' AS='0.105e-6*Wp' PD='Wp+210e-9' PS='Wp+210e-9' M=1
.ends TG_DFSR
